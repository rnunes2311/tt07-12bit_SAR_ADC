VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rnunes2311_12bit_sar_adc
  CLASS BLOCK ;
  FOREIGN tt_um_rnunes2311_12bit_sar_adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.794000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 73.040001 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 88.159996 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 50.680000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.360000 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.360000 ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 63.217499 ;
    ANTENNADIFFAREA 426.674683 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 158.500 5.000 160.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 14.005 217.690 14.175 217.880 ;
        RECT 17.685 217.690 17.855 217.880 ;
        RECT 19.525 217.690 19.695 217.880 ;
        RECT 21.365 217.690 21.535 217.880 ;
        RECT 21.835 217.690 22.005 217.880 ;
        RECT 23.205 217.690 23.375 217.880 ;
        RECT 25.040 217.740 25.160 217.850 ;
        RECT 26.425 217.690 26.595 217.880 ;
        RECT 27.620 217.690 27.790 217.880 ;
        RECT 31.485 217.690 31.655 217.880 ;
        RECT 34.245 217.690 34.415 217.880 ;
        RECT 36.545 217.690 36.715 217.880 ;
        RECT 37.005 217.690 37.175 217.880 ;
        RECT 40.500 217.690 40.670 217.880 ;
        RECT 44.640 217.690 44.810 217.880 ;
        RECT 49.425 217.690 49.595 217.880 ;
        RECT 49.885 217.690 50.055 217.880 ;
        RECT 53.380 217.690 53.550 217.880 ;
        RECT 57.245 217.690 57.415 217.880 ;
        RECT 60.925 217.690 61.095 217.880 ;
        RECT 61.395 217.735 61.555 217.845 ;
        RECT 63.225 217.690 63.395 217.880 ;
        RECT 63.685 217.690 63.855 217.880 ;
        RECT 65.060 217.740 65.180 217.850 ;
        RECT 65.985 217.690 66.155 217.880 ;
        RECT 68.740 217.740 68.860 217.850 ;
        RECT 69.205 217.710 69.375 217.880 ;
        RECT 69.225 217.690 69.375 217.710 ;
        RECT 71.505 217.690 71.675 217.880 ;
        RECT 75.185 217.690 75.355 217.880 ;
        RECT 77.940 217.740 78.060 217.850 ;
        RECT 80.705 217.710 80.875 217.880 ;
        RECT 80.705 217.690 80.855 217.710 ;
        RECT 81.165 217.690 81.335 217.880 ;
        RECT 84.845 217.710 85.015 217.880 ;
        RECT 84.865 217.690 85.015 217.710 ;
        RECT 87.145 217.690 87.315 217.880 ;
        RECT 89.905 217.690 90.075 217.880 ;
        RECT 91.745 217.690 91.915 217.880 ;
        RECT 94.500 217.740 94.620 217.850 ;
        RECT 95.885 217.690 96.055 217.880 ;
        RECT 96.345 217.690 96.515 217.880 ;
        RECT 101.415 217.690 101.585 217.880 ;
        RECT 102.785 217.690 102.955 217.880 ;
        RECT 104.625 217.690 104.795 217.880 ;
        RECT 106.475 217.735 106.635 217.845 ;
        RECT 107.385 217.690 107.555 217.880 ;
        RECT 119.805 217.690 119.975 217.880 ;
        RECT 122.565 217.690 122.735 217.880 ;
        RECT 123.020 217.740 123.140 217.850 ;
        RECT 124.865 217.690 125.035 217.880 ;
        RECT 125.335 217.735 125.495 217.845 ;
        RECT 128.080 217.690 128.250 217.880 ;
        RECT 129.465 217.690 129.635 217.880 ;
        RECT 130.385 217.690 130.555 217.880 ;
        RECT 138.230 217.710 138.400 217.880 ;
        RECT 138.230 217.690 138.340 217.710 ;
        RECT 139.585 217.690 139.755 217.880 ;
        RECT 140.055 217.735 140.215 217.845 ;
        RECT 140.965 217.690 141.135 217.880 ;
        RECT 144.185 217.690 144.355 217.880 ;
        RECT 144.645 217.690 144.815 217.880 ;
        RECT 147.405 217.690 147.575 217.880 ;
        RECT 13.865 216.880 15.235 217.690 ;
        RECT 15.255 217.010 17.995 217.690 ;
        RECT 18.005 217.010 19.835 217.690 ;
        RECT 19.845 217.010 21.675 217.690 ;
        RECT 18.005 216.780 19.350 217.010 ;
        RECT 19.845 216.780 21.190 217.010 ;
        RECT 21.685 216.910 23.055 217.690 ;
        RECT 23.065 216.880 24.895 217.690 ;
        RECT 25.375 216.780 26.725 217.690 ;
        RECT 26.755 216.820 27.185 217.605 ;
        RECT 27.205 217.010 31.105 217.690 ;
        RECT 31.345 217.010 34.085 217.690 ;
        RECT 27.205 216.780 28.135 217.010 ;
        RECT 34.105 216.880 35.475 217.690 ;
        RECT 35.495 216.780 36.845 217.690 ;
        RECT 36.865 217.010 39.605 217.690 ;
        RECT 39.635 216.820 40.065 217.605 ;
        RECT 40.085 217.010 43.985 217.690 ;
        RECT 44.225 217.010 48.125 217.690 ;
        RECT 40.085 216.780 41.015 217.010 ;
        RECT 44.225 216.780 45.155 217.010 ;
        RECT 48.375 216.780 49.725 217.690 ;
        RECT 49.745 217.010 52.485 217.690 ;
        RECT 52.515 216.820 52.945 217.605 ;
        RECT 52.965 217.010 56.865 217.690 ;
        RECT 52.965 216.780 53.895 217.010 ;
        RECT 57.105 216.880 58.475 217.690 ;
        RECT 58.495 217.010 61.235 217.690 ;
        RECT 62.175 216.780 63.525 217.690 ;
        RECT 63.555 216.780 64.905 217.690 ;
        RECT 65.395 216.820 65.825 217.605 ;
        RECT 65.845 217.010 68.585 217.690 ;
        RECT 69.225 216.870 71.155 217.690 ;
        RECT 71.365 216.880 75.035 217.690 ;
        RECT 75.045 217.010 77.785 217.690 ;
        RECT 70.205 216.780 71.155 216.870 ;
        RECT 78.275 216.820 78.705 217.605 ;
        RECT 78.925 216.870 80.855 217.690 ;
        RECT 81.025 216.880 84.695 217.690 ;
        RECT 84.865 216.870 86.795 217.690 ;
        RECT 87.005 217.010 89.745 217.690 ;
        RECT 89.765 216.880 91.135 217.690 ;
        RECT 78.925 216.780 79.875 216.870 ;
        RECT 85.845 216.780 86.795 216.870 ;
        RECT 91.155 216.820 91.585 217.605 ;
        RECT 91.605 216.880 94.355 217.690 ;
        RECT 94.835 216.780 96.185 217.690 ;
        RECT 96.345 217.460 101.250 217.690 ;
        RECT 96.205 216.780 101.250 217.460 ;
        RECT 101.265 216.910 102.635 217.690 ;
        RECT 102.645 216.880 104.015 217.690 ;
        RECT 104.035 216.820 104.465 217.605 ;
        RECT 104.485 217.010 106.315 217.690 ;
        RECT 107.245 217.010 116.855 217.690 ;
        RECT 104.970 216.780 106.315 217.010 ;
        RECT 111.755 216.790 112.685 217.010 ;
        RECT 115.515 216.780 116.855 217.010 ;
        RECT 116.915 216.820 117.345 217.605 ;
        RECT 117.375 217.010 120.115 217.690 ;
        RECT 120.135 217.010 122.875 217.690 ;
        RECT 123.345 217.010 125.175 217.690 ;
        RECT 126.560 217.460 128.250 217.690 ;
        RECT 123.345 216.780 124.690 217.010 ;
        RECT 126.560 216.780 128.395 217.460 ;
        RECT 128.405 216.910 129.775 217.690 ;
        RECT 129.795 216.820 130.225 217.605 ;
        RECT 130.245 216.880 133.915 217.690 ;
        RECT 133.925 217.010 138.340 217.690 ;
        RECT 133.925 216.780 137.855 217.010 ;
        RECT 138.525 216.910 139.895 217.690 ;
        RECT 140.825 217.010 142.655 217.690 ;
        RECT 141.310 216.780 142.655 217.010 ;
        RECT 142.675 216.820 143.105 217.605 ;
        RECT 143.125 216.910 144.495 217.690 ;
        RECT 144.505 217.010 146.335 217.690 ;
        RECT 144.990 216.780 146.335 217.010 ;
        RECT 146.345 216.880 147.715 217.690 ;
      LAYER nwell ;
        RECT 13.670 213.660 147.910 216.490 ;
      LAYER pwell ;
        RECT 13.865 212.460 15.235 213.270 ;
        RECT 15.245 213.140 16.590 213.370 ;
        RECT 17.085 213.140 18.430 213.370 ;
        RECT 18.925 213.140 20.270 213.370 ;
        RECT 25.585 213.280 26.535 213.370 ;
        RECT 15.245 212.460 17.075 213.140 ;
        RECT 17.085 212.460 18.915 213.140 ;
        RECT 18.925 212.460 20.755 213.140 ;
        RECT 20.765 212.460 24.435 213.270 ;
        RECT 24.605 212.460 26.535 213.280 ;
        RECT 26.755 212.545 27.185 213.330 ;
        RECT 27.205 212.460 29.035 213.270 ;
        RECT 33.555 213.140 34.485 213.360 ;
        RECT 37.205 213.140 39.415 213.370 ;
        RECT 29.045 212.460 39.415 213.140 ;
        RECT 39.625 212.690 41.460 213.370 ;
        RECT 46.435 213.140 47.365 213.360 ;
        RECT 50.195 213.140 51.115 213.370 ;
        RECT 39.770 212.460 41.460 212.690 ;
        RECT 41.925 212.460 51.115 213.140 ;
        RECT 51.125 212.460 52.495 213.270 ;
        RECT 52.515 212.545 52.945 213.330 ;
        RECT 57.475 213.140 58.405 213.360 ;
        RECT 61.235 213.140 62.155 213.370 ;
        RECT 52.965 212.460 62.155 213.140 ;
        RECT 62.165 213.140 63.095 213.370 ;
        RECT 71.275 213.140 72.205 213.360 ;
        RECT 75.035 213.140 76.375 213.370 ;
        RECT 62.165 212.460 66.065 213.140 ;
        RECT 66.765 212.460 76.375 213.140 ;
        RECT 76.435 212.460 77.785 213.370 ;
        RECT 78.275 212.545 78.705 213.330 ;
        RECT 78.765 213.140 80.105 213.370 ;
        RECT 82.935 213.140 83.865 213.360 ;
        RECT 92.895 213.140 93.825 213.360 ;
        RECT 96.655 213.140 97.575 213.370 ;
        RECT 98.725 213.280 99.675 213.370 ;
        RECT 78.765 212.460 88.375 213.140 ;
        RECT 88.385 212.460 97.575 213.140 ;
        RECT 97.745 212.460 99.675 213.280 ;
        RECT 99.885 213.140 100.815 213.370 ;
        RECT 99.885 212.460 103.785 213.140 ;
        RECT 104.035 212.545 104.465 213.330 ;
        RECT 104.495 212.460 107.225 213.370 ;
        RECT 107.245 212.460 109.075 213.140 ;
        RECT 109.085 212.460 110.915 213.270 ;
        RECT 110.925 213.140 111.855 213.370 ;
        RECT 110.925 212.460 114.825 213.140 ;
        RECT 115.995 212.460 117.345 213.370 ;
        RECT 117.495 212.460 123.335 213.370 ;
        RECT 123.800 212.690 125.635 213.370 ;
        RECT 123.800 212.460 125.490 212.690 ;
        RECT 126.115 212.460 128.845 213.370 ;
        RECT 129.795 212.545 130.225 213.330 ;
        RECT 134.755 213.140 135.685 213.360 ;
        RECT 138.515 213.140 139.435 213.370 ;
        RECT 130.245 212.460 139.435 213.140 ;
        RECT 139.445 213.140 140.790 213.370 ;
        RECT 139.445 212.460 141.275 213.140 ;
        RECT 141.285 212.460 142.655 213.240 ;
        RECT 143.150 213.140 144.495 213.370 ;
        RECT 144.990 213.140 146.335 213.370 ;
        RECT 142.665 212.460 144.495 213.140 ;
        RECT 144.505 212.460 146.335 213.140 ;
        RECT 146.345 212.460 147.715 213.270 ;
        RECT 14.005 212.250 14.175 212.460 ;
        RECT 16.765 212.250 16.935 212.460 ;
        RECT 18.605 212.250 18.775 212.460 ;
        RECT 19.065 212.250 19.235 212.440 ;
        RECT 20.445 212.270 20.615 212.460 ;
        RECT 20.905 212.270 21.075 212.460 ;
        RECT 24.605 212.440 24.755 212.460 ;
        RECT 24.585 212.270 24.755 212.440 ;
        RECT 27.345 212.270 27.515 212.460 ;
        RECT 29.185 212.270 29.355 212.460 ;
        RECT 29.645 212.250 29.815 212.440 ;
        RECT 31.760 212.250 31.930 212.440 ;
        RECT 35.630 212.250 35.800 212.440 ;
        RECT 38.855 212.295 39.015 212.405 ;
        RECT 39.770 212.270 39.940 212.460 ;
        RECT 40.220 212.300 40.340 212.410 ;
        RECT 40.660 212.270 40.830 212.440 ;
        RECT 42.065 212.270 42.235 212.460 ;
        RECT 40.720 212.250 40.830 212.270 ;
        RECT 47.585 212.250 47.755 212.440 ;
        RECT 49.885 212.270 50.055 212.440 ;
        RECT 50.355 212.295 50.515 212.405 ;
        RECT 51.265 212.270 51.435 212.460 ;
        RECT 49.885 212.250 50.035 212.270 ;
        RECT 52.190 212.250 52.360 212.440 ;
        RECT 52.640 212.300 52.760 212.410 ;
        RECT 53.105 212.270 53.275 212.460 ;
        RECT 54.485 212.250 54.655 212.440 ;
        RECT 55.220 212.250 55.390 212.440 ;
        RECT 60.005 212.250 60.175 212.440 ;
        RECT 62.580 212.270 62.750 212.460 ;
        RECT 63.870 212.250 64.040 212.440 ;
        RECT 64.615 212.295 64.775 212.405 ;
        RECT 65.985 212.250 66.155 212.440 ;
        RECT 66.440 212.300 66.560 212.410 ;
        RECT 66.905 212.270 67.075 212.460 ;
        RECT 76.565 212.440 76.735 212.460 ;
        RECT 68.740 212.300 68.860 212.410 ;
        RECT 69.480 212.250 69.650 212.440 ;
        RECT 74.270 212.250 74.440 212.440 ;
        RECT 74.735 212.295 74.895 212.405 ;
        RECT 76.565 212.270 76.740 212.440 ;
        RECT 77.020 212.300 77.140 212.410 ;
        RECT 77.940 212.300 78.060 212.410 ;
        RECT 76.570 212.250 76.740 212.270 ;
        RECT 80.890 212.250 81.060 212.440 ;
        RECT 81.625 212.250 81.795 212.440 ;
        RECT 84.385 212.250 84.555 212.440 ;
        RECT 84.840 212.300 84.960 212.410 ;
        RECT 88.065 212.270 88.235 212.460 ;
        RECT 88.525 212.270 88.695 212.460 ;
        RECT 97.745 212.440 97.895 212.460 ;
        RECT 88.710 212.250 88.880 212.440 ;
        RECT 89.440 212.250 89.610 212.440 ;
        RECT 90.820 212.300 90.940 212.410 ;
        RECT 91.745 212.250 91.915 212.440 ;
        RECT 97.725 212.250 97.895 212.440 ;
        RECT 98.180 212.300 98.300 212.410 ;
        RECT 98.645 212.250 98.815 212.440 ;
        RECT 100.300 212.270 100.470 212.460 ;
        RECT 104.625 212.270 104.795 212.460 ;
        RECT 107.845 212.250 108.015 212.440 ;
        RECT 108.765 212.270 108.935 212.460 ;
        RECT 109.225 212.270 109.395 212.460 ;
        RECT 111.340 212.270 111.510 212.460 ;
        RECT 115.215 212.305 115.375 212.415 ;
        RECT 116.125 212.270 116.295 212.460 ;
        RECT 118.885 212.250 119.055 212.440 ;
        RECT 122.100 212.250 122.270 212.440 ;
        RECT 123.025 212.270 123.195 212.460 ;
        RECT 123.485 212.250 123.655 212.440 ;
        RECT 123.945 212.250 124.115 212.440 ;
        RECT 125.320 212.270 125.490 212.460 ;
        RECT 125.780 212.300 125.900 212.410 ;
        RECT 126.245 212.270 126.415 212.460 ;
        RECT 129.015 212.305 129.175 212.415 ;
        RECT 130.385 212.270 130.555 212.460 ;
        RECT 133.420 212.250 133.590 212.440 ;
        RECT 137.285 212.250 137.455 212.440 ;
        RECT 140.965 212.250 141.135 212.460 ;
        RECT 142.335 212.270 142.505 212.460 ;
        RECT 142.805 212.270 142.975 212.460 ;
        RECT 143.265 212.250 143.435 212.440 ;
        RECT 144.645 212.250 144.815 212.460 ;
        RECT 147.405 212.250 147.575 212.460 ;
        RECT 13.865 211.440 15.235 212.250 ;
        RECT 15.245 211.570 17.075 212.250 ;
        RECT 17.085 211.570 18.915 212.250 ;
        RECT 18.925 211.570 29.295 212.250 ;
        RECT 15.245 211.340 16.590 211.570 ;
        RECT 17.085 211.340 18.430 211.570 ;
        RECT 23.435 211.350 24.365 211.570 ;
        RECT 27.085 211.340 29.295 211.570 ;
        RECT 29.505 211.440 31.335 212.250 ;
        RECT 31.345 211.570 35.245 212.250 ;
        RECT 31.345 211.340 32.275 211.570 ;
        RECT 35.485 211.340 38.405 212.250 ;
        RECT 39.635 211.380 40.065 212.165 ;
        RECT 40.720 211.570 45.135 212.250 ;
        RECT 45.155 211.570 47.895 212.250 ;
        RECT 41.205 211.340 45.135 211.570 ;
        RECT 48.105 211.430 50.035 212.250 ;
        RECT 48.105 211.340 49.055 211.430 ;
        RECT 51.125 211.340 52.475 212.250 ;
        RECT 52.965 211.570 54.795 212.250 ;
        RECT 54.805 211.570 58.705 212.250 ;
        RECT 52.965 211.340 54.310 211.570 ;
        RECT 54.805 211.340 55.735 211.570 ;
        RECT 58.955 211.340 60.305 212.250 ;
        RECT 60.555 211.570 64.455 212.250 ;
        RECT 63.525 211.340 64.455 211.570 ;
        RECT 65.395 211.380 65.825 212.165 ;
        RECT 65.845 211.440 68.595 212.250 ;
        RECT 69.065 211.570 72.965 212.250 ;
        RECT 69.065 211.340 69.995 211.570 ;
        RECT 73.205 211.340 74.555 212.250 ;
        RECT 75.505 211.340 76.855 212.250 ;
        RECT 77.575 211.570 81.475 212.250 ;
        RECT 81.485 211.570 83.315 212.250 ;
        RECT 80.545 211.340 81.475 211.570 ;
        RECT 83.335 211.340 84.685 212.250 ;
        RECT 85.395 211.570 89.295 212.250 ;
        RECT 88.365 211.340 89.295 211.570 ;
        RECT 89.325 211.340 90.675 212.250 ;
        RECT 91.155 211.380 91.585 212.165 ;
        RECT 91.605 211.340 96.155 212.250 ;
        RECT 96.205 211.570 98.035 212.250 ;
        RECT 98.505 211.570 107.695 212.250 ;
        RECT 107.705 211.570 116.810 212.250 ;
        RECT 103.015 211.350 103.945 211.570 ;
        RECT 106.775 211.340 107.695 211.570 ;
        RECT 116.915 211.380 117.345 212.165 ;
        RECT 117.365 211.570 119.195 212.250 ;
        RECT 119.495 211.340 122.415 212.250 ;
        RECT 122.435 211.340 123.785 212.250 ;
        RECT 123.805 211.570 132.995 212.250 ;
        RECT 128.315 211.350 129.245 211.570 ;
        RECT 132.075 211.340 132.995 211.570 ;
        RECT 133.005 211.570 136.905 212.250 ;
        RECT 133.005 211.340 133.935 211.570 ;
        RECT 137.145 211.440 140.815 212.250 ;
        RECT 140.825 211.570 142.655 212.250 ;
        RECT 141.310 211.340 142.655 211.570 ;
        RECT 142.675 211.380 143.105 212.165 ;
        RECT 143.125 211.440 144.495 212.250 ;
        RECT 144.505 211.570 146.335 212.250 ;
        RECT 144.990 211.340 146.335 211.570 ;
        RECT 146.345 211.440 147.715 212.250 ;
      LAYER nwell ;
        RECT 13.670 208.220 147.910 211.050 ;
      LAYER pwell ;
        RECT 13.865 207.020 15.235 207.830 ;
        RECT 15.245 207.700 16.590 207.930 ;
        RECT 17.085 207.700 18.430 207.930 ;
        RECT 15.245 207.020 17.075 207.700 ;
        RECT 17.085 207.020 18.915 207.700 ;
        RECT 18.925 207.020 22.595 207.830 ;
        RECT 22.605 207.020 23.975 207.830 ;
        RECT 24.215 207.250 26.605 207.930 ;
        RECT 24.215 207.020 26.595 207.250 ;
        RECT 26.755 207.105 27.185 207.890 ;
        RECT 27.205 207.700 28.135 207.930 ;
        RECT 27.205 207.020 31.105 207.700 ;
        RECT 31.345 207.020 34.265 207.930 ;
        RECT 34.695 207.250 37.085 207.930 ;
        RECT 34.705 207.020 37.085 207.250 ;
        RECT 37.345 207.020 38.695 207.930 ;
        RECT 38.705 207.700 39.635 207.930 ;
        RECT 38.705 207.020 42.605 207.700 ;
        RECT 42.855 207.020 44.205 207.930 ;
        RECT 44.235 207.020 46.965 207.930 ;
        RECT 46.985 207.730 47.930 207.930 ;
        RECT 49.265 207.730 50.195 207.930 ;
        RECT 46.985 207.250 50.195 207.730 ;
        RECT 50.690 207.700 52.035 207.930 ;
        RECT 46.985 207.050 50.055 207.250 ;
        RECT 46.985 207.020 47.930 207.050 ;
        RECT 14.005 206.810 14.175 207.020 ;
        RECT 16.765 206.810 16.935 207.020 ;
        RECT 18.605 206.810 18.775 207.020 ;
        RECT 19.065 206.830 19.235 207.020 ;
        RECT 19.985 206.810 20.155 207.000 ;
        RECT 20.445 206.810 20.615 207.000 ;
        RECT 22.745 206.830 22.915 207.020 ;
        RECT 24.120 206.860 24.240 206.970 ;
        RECT 25.500 206.810 25.670 207.000 ;
        RECT 25.965 206.830 26.135 207.000 ;
        RECT 26.425 206.830 26.595 207.020 ;
        RECT 27.620 206.830 27.790 207.020 ;
        RECT 28.260 206.860 28.380 206.970 ;
        RECT 25.985 206.810 26.135 206.830 ;
        RECT 13.865 206.000 15.235 206.810 ;
        RECT 15.245 206.130 17.075 206.810 ;
        RECT 17.085 206.130 18.915 206.810 ;
        RECT 15.245 205.900 16.590 206.130 ;
        RECT 17.085 205.900 18.430 206.130 ;
        RECT 18.925 206.030 20.295 206.810 ;
        RECT 20.305 206.000 23.975 206.810 ;
        RECT 24.465 205.900 25.815 206.810 ;
        RECT 25.985 205.990 27.915 206.810 ;
        RECT 28.725 206.780 28.895 207.000 ;
        RECT 31.490 206.830 31.660 207.020 ;
        RECT 32.870 206.810 33.040 207.000 ;
        RECT 33.325 206.810 33.495 207.000 ;
        RECT 34.705 206.830 34.875 207.020 ;
        RECT 36.090 206.810 36.260 207.000 ;
        RECT 36.545 206.810 36.715 207.000 ;
        RECT 37.460 206.830 37.630 207.020 ;
        RECT 39.120 206.830 39.290 207.020 ;
        RECT 42.985 207.000 43.155 207.020 ;
        RECT 39.305 206.810 39.475 207.000 ;
        RECT 42.525 206.810 42.695 207.000 ;
        RECT 42.985 206.830 43.160 207.000 ;
        RECT 44.365 206.830 44.535 207.020 ;
        RECT 46.200 206.860 46.320 206.970 ;
        RECT 42.990 206.810 43.160 206.830 ;
        RECT 48.965 206.810 49.135 207.000 ;
        RECT 49.435 206.855 49.595 206.965 ;
        RECT 49.885 206.830 50.055 207.050 ;
        RECT 50.205 207.020 52.035 207.700 ;
        RECT 52.515 207.105 52.945 207.890 ;
        RECT 52.995 207.020 55.715 207.930 ;
        RECT 55.925 207.840 56.875 207.930 ;
        RECT 55.925 207.020 57.855 207.840 ;
        RECT 58.985 207.700 60.325 207.930 ;
        RECT 63.155 207.700 64.085 207.920 ;
        RECT 58.985 207.020 68.595 207.700 ;
        RECT 69.555 207.020 72.275 207.930 ;
        RECT 72.285 207.020 75.205 207.930 ;
        RECT 75.505 207.020 77.335 207.930 ;
        RECT 78.275 207.105 78.705 207.890 ;
        RECT 79.645 207.020 83.315 207.930 ;
        RECT 84.275 207.020 86.995 207.930 ;
        RECT 87.005 207.020 90.675 207.930 ;
        RECT 91.605 207.700 92.535 207.930 ;
        RECT 95.285 207.700 96.215 207.930 ;
        RECT 91.605 207.020 95.275 207.700 ;
        RECT 95.285 207.020 98.955 207.700 ;
        RECT 98.965 207.020 101.885 207.930 ;
        RECT 102.185 207.020 104.015 207.700 ;
        RECT 104.035 207.105 104.465 207.890 ;
        RECT 104.485 207.730 105.415 207.930 ;
        RECT 106.750 207.730 107.695 207.930 ;
        RECT 104.485 207.250 107.695 207.730 ;
        RECT 112.215 207.700 113.145 207.920 ;
        RECT 115.975 207.700 116.895 207.930 ;
        RECT 104.625 207.050 107.695 207.250 ;
        RECT 50.345 207.000 50.515 207.020 ;
        RECT 50.340 206.830 50.515 207.000 ;
        RECT 51.720 206.860 51.840 206.970 ;
        RECT 52.180 206.860 52.300 206.970 ;
        RECT 50.340 206.810 50.510 206.830 ;
        RECT 54.020 206.810 54.190 207.000 ;
        RECT 54.490 206.810 54.660 207.000 ;
        RECT 55.405 206.830 55.575 207.020 ;
        RECT 57.705 207.000 57.855 207.020 ;
        RECT 57.705 206.830 57.875 207.000 ;
        RECT 58.175 206.865 58.335 206.975 ;
        RECT 60.925 206.810 61.095 207.000 ;
        RECT 61.380 206.860 61.500 206.970 ;
        RECT 61.845 206.830 62.015 207.000 ;
        RECT 61.865 206.810 62.015 206.830 ;
        RECT 64.140 206.810 64.310 207.000 ;
        RECT 66.260 206.810 66.430 207.000 ;
        RECT 68.285 206.830 68.455 207.020 ;
        RECT 68.755 206.865 68.915 206.975 ;
        RECT 71.050 206.810 71.220 207.000 ;
        RECT 71.965 206.830 72.135 207.020 ;
        RECT 72.430 206.830 72.600 207.020 ;
        RECT 73.805 206.810 73.975 207.000 ;
        RECT 75.650 206.830 75.820 207.020 ;
        RECT 77.495 206.865 77.655 206.975 ;
        RECT 78.875 206.865 79.035 206.975 ;
        RECT 79.790 206.830 79.960 207.020 ;
        RECT 83.005 206.810 83.175 207.000 ;
        RECT 83.475 206.865 83.635 206.975 ;
        RECT 85.765 206.810 85.935 207.000 ;
        RECT 86.220 206.810 86.390 207.000 ;
        RECT 86.685 206.830 86.855 207.020 ;
        RECT 87.150 206.830 87.320 207.020 ;
        RECT 87.615 206.855 87.775 206.965 ;
        RECT 90.825 206.810 90.995 207.000 ;
        RECT 92.665 206.810 92.835 207.000 ;
        RECT 93.125 206.810 93.295 207.000 ;
        RECT 94.965 206.830 95.135 207.020 ;
        RECT 95.890 206.810 96.060 207.000 ;
        RECT 96.620 206.810 96.790 207.000 ;
        RECT 98.645 206.830 98.815 207.020 ;
        RECT 99.110 206.830 99.280 207.020 ;
        RECT 100.490 206.810 100.660 207.000 ;
        RECT 102.325 206.830 102.495 207.020 ;
        RECT 103.705 206.810 103.875 207.000 ;
        RECT 104.625 206.830 104.795 207.050 ;
        RECT 106.750 207.020 107.695 207.050 ;
        RECT 107.705 207.020 116.895 207.700 ;
        RECT 117.100 207.020 120.575 207.930 ;
        RECT 125.095 207.700 126.025 207.920 ;
        RECT 128.855 207.700 129.775 207.930 ;
        RECT 120.585 207.020 129.775 207.700 ;
        RECT 129.795 207.105 130.225 207.890 ;
        RECT 134.755 207.700 135.685 207.920 ;
        RECT 138.515 207.700 139.435 207.930 ;
        RECT 130.245 207.020 139.435 207.700 ;
        RECT 139.445 207.020 140.815 207.830 ;
        RECT 141.310 207.700 142.655 207.930 ;
        RECT 143.150 207.700 144.495 207.930 ;
        RECT 144.990 207.700 146.335 207.930 ;
        RECT 140.825 207.020 142.655 207.700 ;
        RECT 142.665 207.020 144.495 207.700 ;
        RECT 144.505 207.020 146.335 207.700 ;
        RECT 146.345 207.020 147.715 207.830 ;
        RECT 106.460 206.860 106.580 206.970 ;
        RECT 106.925 206.810 107.095 207.000 ;
        RECT 107.845 206.830 108.015 207.020 ;
        RECT 109.690 206.810 109.860 207.000 ;
        RECT 30.850 206.780 31.795 206.810 ;
        RECT 28.725 206.580 31.795 206.780 ;
        RECT 26.965 205.900 27.915 205.990 ;
        RECT 28.585 206.100 31.795 206.580 ;
        RECT 28.585 205.900 29.515 206.100 ;
        RECT 30.850 205.900 31.795 206.100 ;
        RECT 31.805 205.900 33.155 206.810 ;
        RECT 33.185 206.000 35.015 206.810 ;
        RECT 35.025 205.900 36.375 206.810 ;
        RECT 36.415 205.900 37.765 206.810 ;
        RECT 37.785 206.130 39.615 206.810 ;
        RECT 39.635 205.940 40.065 206.725 ;
        RECT 40.115 205.900 42.835 206.810 ;
        RECT 42.845 205.900 45.765 206.810 ;
        RECT 46.755 206.580 49.135 206.810 ;
        RECT 46.755 205.900 49.145 206.580 ;
        RECT 50.225 205.900 51.575 206.810 ;
        RECT 52.500 206.580 54.190 206.810 ;
        RECT 52.500 205.900 54.335 206.580 ;
        RECT 54.345 205.900 58.000 206.810 ;
        RECT 58.025 205.900 61.235 206.810 ;
        RECT 61.865 205.990 63.795 206.810 ;
        RECT 62.845 205.900 63.795 205.990 ;
        RECT 64.025 205.900 65.375 206.810 ;
        RECT 65.395 205.940 65.825 206.725 ;
        RECT 65.845 206.130 69.745 206.810 ;
        RECT 65.845 205.900 66.775 206.130 ;
        RECT 69.985 205.900 71.335 206.810 ;
        RECT 71.395 205.900 74.115 206.810 ;
        RECT 74.210 206.130 83.315 206.810 ;
        RECT 83.325 206.130 86.075 206.810 ;
        RECT 83.325 205.900 84.255 206.130 ;
        RECT 86.105 205.900 87.455 206.810 ;
        RECT 88.385 206.130 91.135 206.810 ;
        RECT 88.385 205.900 89.315 206.130 ;
        RECT 91.155 205.940 91.585 206.725 ;
        RECT 91.615 205.900 92.965 206.810 ;
        RECT 92.985 206.000 94.815 206.810 ;
        RECT 94.825 205.900 96.175 206.810 ;
        RECT 96.205 206.130 100.105 206.810 ;
        RECT 96.205 205.900 97.135 206.130 ;
        RECT 100.345 205.900 103.265 206.810 ;
        RECT 103.705 206.580 106.085 206.810 ;
        RECT 103.695 205.900 106.085 206.580 ;
        RECT 106.785 206.130 109.535 206.810 ;
        RECT 108.605 205.900 109.535 206.130 ;
        RECT 109.545 205.900 113.215 206.810 ;
        RECT 113.225 206.780 114.170 206.810 ;
        RECT 116.125 206.780 116.295 207.000 ;
        RECT 116.580 206.860 116.700 206.970 ;
        RECT 117.510 206.780 117.680 207.000 ;
        RECT 120.260 206.830 120.430 207.020 ;
        RECT 120.725 206.830 120.895 207.020 ;
        RECT 120.085 206.780 121.035 206.810 ;
        RECT 113.225 206.580 116.295 206.780 ;
        RECT 113.225 206.100 116.435 206.580 ;
        RECT 113.225 205.900 114.170 206.100 ;
        RECT 115.505 205.900 116.435 206.100 ;
        RECT 116.915 205.940 117.345 206.725 ;
        RECT 117.365 206.100 121.035 206.780 ;
        RECT 120.085 205.900 121.035 206.100 ;
        RECT 121.045 206.780 121.990 206.810 ;
        RECT 123.945 206.780 124.115 207.000 ;
        RECT 121.045 206.580 124.115 206.780 ;
        RECT 124.410 206.810 124.580 207.000 ;
        RECT 127.625 206.810 127.795 207.000 ;
        RECT 129.920 206.810 130.090 207.000 ;
        RECT 130.385 206.830 130.555 207.020 ;
        RECT 131.300 206.810 131.470 207.000 ;
        RECT 131.775 206.855 131.935 206.965 ;
        RECT 132.685 206.810 132.855 207.000 ;
        RECT 137.745 206.810 137.915 207.000 ;
        RECT 138.205 206.810 138.375 207.000 ;
        RECT 139.585 206.830 139.755 207.020 ;
        RECT 140.965 206.810 141.135 207.020 ;
        RECT 142.805 206.830 142.975 207.020 ;
        RECT 143.265 206.810 143.435 207.000 ;
        RECT 144.645 206.810 144.815 207.020 ;
        RECT 147.405 206.810 147.575 207.020 ;
        RECT 124.410 206.580 127.465 206.810 ;
        RECT 121.045 206.100 124.255 206.580 ;
        RECT 121.045 205.900 121.990 206.100 ;
        RECT 123.325 205.900 124.255 206.100 ;
        RECT 124.265 205.900 127.465 206.580 ;
        RECT 127.495 205.900 128.845 206.810 ;
        RECT 128.885 205.900 130.235 206.810 ;
        RECT 130.265 205.900 131.615 206.810 ;
        RECT 132.545 206.130 134.375 206.810 ;
        RECT 133.030 205.900 134.375 206.130 ;
        RECT 134.480 206.130 137.945 206.810 ;
        RECT 134.480 205.900 135.400 206.130 ;
        RECT 138.065 206.000 140.815 206.810 ;
        RECT 140.825 206.130 142.655 206.810 ;
        RECT 141.310 205.900 142.655 206.130 ;
        RECT 142.675 205.940 143.105 206.725 ;
        RECT 143.125 206.000 144.495 206.810 ;
        RECT 144.505 206.130 146.335 206.810 ;
        RECT 144.990 205.900 146.335 206.130 ;
        RECT 146.345 206.000 147.715 206.810 ;
      LAYER nwell ;
        RECT 13.670 202.780 147.910 205.610 ;
      LAYER pwell ;
        RECT 13.865 201.580 15.235 202.390 ;
        RECT 15.245 202.260 16.590 202.490 ;
        RECT 22.055 202.260 22.985 202.480 ;
        RECT 25.815 202.260 26.735 202.490 ;
        RECT 15.245 201.580 17.075 202.260 ;
        RECT 17.545 201.580 26.735 202.260 ;
        RECT 26.755 201.665 27.185 202.450 ;
        RECT 27.205 202.260 28.135 202.490 ;
        RECT 27.205 201.580 31.105 202.260 ;
        RECT 31.375 201.580 34.095 202.490 ;
        RECT 34.190 201.580 43.295 202.260 ;
        RECT 43.315 201.580 46.055 202.260 ;
        RECT 46.525 201.580 48.715 202.490 ;
        RECT 48.835 201.580 50.185 202.490 ;
        RECT 50.205 201.580 51.555 202.490 ;
        RECT 52.515 201.665 52.945 202.450 ;
        RECT 53.425 201.580 55.255 202.260 ;
        RECT 55.325 201.580 57.095 202.490 ;
        RECT 57.300 201.580 60.775 202.490 ;
        RECT 69.985 202.290 70.930 202.490 ;
        RECT 72.265 202.290 73.195 202.490 ;
        RECT 74.540 202.290 75.495 202.490 ;
        RECT 60.785 201.580 69.890 202.260 ;
        RECT 69.985 201.810 73.195 202.290 ;
        RECT 69.985 201.610 73.055 201.810 ;
        RECT 73.215 201.610 75.495 202.290 ;
        RECT 69.985 201.580 70.930 201.610 ;
        RECT 14.005 201.370 14.175 201.580 ;
        RECT 16.765 201.370 16.935 201.580 ;
        RECT 17.220 201.420 17.340 201.530 ;
        RECT 17.685 201.390 17.855 201.580 ;
        RECT 18.605 201.370 18.775 201.560 ;
        RECT 19.060 201.420 19.180 201.530 ;
        RECT 19.525 201.370 19.695 201.560 ;
        RECT 27.620 201.390 27.790 201.580 ;
        RECT 30.100 201.420 30.220 201.530 ;
        RECT 30.565 201.390 30.735 201.560 ;
        RECT 32.865 201.390 33.035 201.560 ;
        RECT 33.785 201.390 33.955 201.580 ;
        RECT 30.585 201.370 30.735 201.390 ;
        RECT 32.870 201.370 33.035 201.390 ;
        RECT 38.380 201.370 38.550 201.560 ;
        RECT 38.855 201.415 39.015 201.525 ;
        RECT 42.985 201.390 43.155 201.580 ;
        RECT 43.440 201.370 43.610 201.560 ;
        RECT 45.745 201.390 45.915 201.580 ;
        RECT 46.210 201.530 46.380 201.560 ;
        RECT 46.200 201.420 46.380 201.530 ;
        RECT 45.745 201.370 45.910 201.390 ;
        RECT 46.210 201.370 46.380 201.420 ;
        RECT 46.670 201.390 46.840 201.580 ;
        RECT 47.575 201.370 47.745 201.560 ;
        RECT 49.885 201.390 50.055 201.580 ;
        RECT 50.350 201.390 50.520 201.580 ;
        RECT 50.805 201.370 50.975 201.560 ;
        RECT 51.735 201.425 51.895 201.535 ;
        RECT 52.185 201.370 52.355 201.560 ;
        RECT 53.100 201.420 53.220 201.530 ;
        RECT 53.565 201.390 53.735 201.580 ;
        RECT 55.400 201.370 55.570 201.560 ;
        RECT 55.865 201.390 56.035 201.560 ;
        RECT 56.780 201.390 56.950 201.580 ;
        RECT 55.870 201.370 56.035 201.390 ;
        RECT 58.170 201.370 58.340 201.560 ;
        RECT 60.460 201.390 60.630 201.580 ;
        RECT 60.925 201.390 61.095 201.580 ;
        RECT 61.845 201.370 62.015 201.560 ;
        RECT 64.615 201.415 64.775 201.525 ;
        RECT 65.985 201.370 66.155 201.560 ;
        RECT 71.045 201.370 71.215 201.560 ;
        RECT 13.865 200.560 15.235 201.370 ;
        RECT 15.245 200.690 17.075 201.370 ;
        RECT 17.085 200.690 18.915 201.370 ;
        RECT 19.385 200.690 29.755 201.370 ;
        RECT 15.245 200.460 16.590 200.690 ;
        RECT 17.085 200.460 18.430 200.690 ;
        RECT 23.895 200.470 24.825 200.690 ;
        RECT 27.545 200.460 29.755 200.690 ;
        RECT 30.585 200.550 32.515 201.370 ;
        RECT 32.870 200.690 34.705 201.370 ;
        RECT 31.565 200.460 32.515 200.550 ;
        RECT 33.775 200.460 34.705 200.690 ;
        RECT 35.040 200.460 38.695 201.370 ;
        RECT 39.635 200.500 40.065 201.285 ;
        RECT 40.100 200.460 43.755 201.370 ;
        RECT 44.075 200.690 45.910 201.370 ;
        RECT 44.075 200.460 45.005 200.690 ;
        RECT 46.065 200.460 47.415 201.370 ;
        RECT 47.445 200.460 50.655 201.370 ;
        RECT 50.675 200.460 52.025 201.370 ;
        RECT 52.055 200.460 53.405 201.370 ;
        RECT 54.365 200.460 55.715 201.370 ;
        RECT 55.870 200.690 57.705 201.370 ;
        RECT 56.775 200.460 57.705 200.690 ;
        RECT 58.025 200.460 61.680 201.370 ;
        RECT 61.715 200.460 64.445 201.370 ;
        RECT 65.395 200.500 65.825 201.285 ;
        RECT 65.855 200.460 68.585 201.370 ;
        RECT 68.835 201.140 71.215 201.370 ;
        RECT 71.500 201.340 71.670 201.560 ;
        RECT 72.885 201.390 73.055 201.610 ;
        RECT 73.340 201.390 73.510 201.610 ;
        RECT 74.540 201.580 75.495 201.610 ;
        RECT 75.505 201.580 77.335 202.490 ;
        RECT 78.275 201.665 78.705 202.450 ;
        RECT 79.385 202.260 83.315 202.490 ;
        RECT 78.900 201.580 83.315 202.260 ;
        RECT 83.345 201.580 84.695 202.490 ;
        RECT 84.715 201.580 86.065 202.490 ;
        RECT 87.005 201.580 88.835 202.490 ;
        RECT 88.845 201.580 90.195 202.490 ;
        RECT 90.245 201.580 91.595 202.490 ;
        RECT 92.065 201.580 93.415 202.490 ;
        RECT 93.445 201.580 94.795 202.490 ;
        RECT 94.825 201.580 98.035 202.490 ;
        RECT 98.045 201.580 101.255 202.490 ;
        RECT 102.205 201.580 103.555 202.490 ;
        RECT 104.035 201.665 104.465 202.450 ;
        RECT 104.485 202.260 105.415 202.490 ;
        RECT 104.485 201.580 108.385 202.260 ;
        RECT 108.635 201.580 109.985 202.490 ;
        RECT 110.005 201.580 112.925 202.490 ;
        RECT 113.245 201.580 114.595 202.490 ;
        RECT 114.605 201.580 117.815 202.490 ;
        RECT 118.285 202.260 119.205 202.490 ;
        RECT 122.035 202.260 122.965 202.480 ;
        RECT 127.685 202.400 128.635 202.490 ;
        RECT 118.285 201.580 127.475 202.260 ;
        RECT 127.685 201.580 129.615 202.400 ;
        RECT 129.795 201.665 130.225 202.450 ;
        RECT 130.245 202.260 131.165 202.490 ;
        RECT 133.995 202.260 134.925 202.480 ;
        RECT 130.245 201.580 139.435 202.260 ;
        RECT 139.455 201.580 140.805 202.490 ;
        RECT 141.285 201.580 142.655 202.360 ;
        RECT 143.150 202.260 144.495 202.490 ;
        RECT 144.990 202.260 146.335 202.490 ;
        RECT 142.665 201.580 144.495 202.260 ;
        RECT 144.505 201.580 146.335 202.260 ;
        RECT 146.345 201.580 147.715 202.390 ;
        RECT 73.815 201.415 73.975 201.525 ;
        RECT 74.715 201.370 74.885 201.560 ;
        RECT 75.650 201.390 75.820 201.580 ;
        RECT 78.900 201.560 79.010 201.580 ;
        RECT 77.495 201.425 77.655 201.535 ;
        RECT 77.950 201.370 78.120 201.560 ;
        RECT 78.840 201.390 79.010 201.560 ;
        RECT 81.160 201.420 81.280 201.530 ;
        RECT 81.620 201.390 81.790 201.560 ;
        RECT 83.460 201.390 83.630 201.580 ;
        RECT 81.655 201.370 81.790 201.390 ;
        RECT 85.310 201.370 85.480 201.560 ;
        RECT 85.765 201.390 85.935 201.580 ;
        RECT 86.235 201.425 86.395 201.535 ;
        RECT 88.520 201.390 88.690 201.580 ;
        RECT 89.910 201.560 90.080 201.580 ;
        RECT 89.900 201.390 90.080 201.560 ;
        RECT 90.360 201.525 90.530 201.580 ;
        RECT 90.360 201.415 90.535 201.525 ;
        RECT 91.740 201.420 91.860 201.530 ;
        RECT 90.360 201.390 90.530 201.415 ;
        RECT 93.130 201.390 93.300 201.580 ;
        RECT 94.510 201.560 94.680 201.580 ;
        RECT 94.505 201.390 94.680 201.560 ;
        RECT 94.955 201.560 95.125 201.580 ;
        RECT 94.955 201.390 95.135 201.560 ;
        RECT 96.800 201.420 96.920 201.530 ;
        RECT 89.900 201.370 90.070 201.390 ;
        RECT 94.505 201.370 94.675 201.390 ;
        RECT 94.965 201.370 95.135 201.390 ;
        RECT 97.265 201.370 97.435 201.560 ;
        RECT 98.175 201.390 98.345 201.580 ;
        RECT 100.485 201.370 100.655 201.560 ;
        RECT 101.415 201.425 101.575 201.535 ;
        RECT 102.320 201.390 102.490 201.580 ;
        RECT 102.790 201.370 102.960 201.560 ;
        RECT 103.700 201.420 103.820 201.530 ;
        RECT 104.170 201.370 104.340 201.560 ;
        RECT 104.625 201.370 104.795 201.560 ;
        RECT 104.900 201.390 105.070 201.580 ;
        RECT 107.845 201.370 108.015 201.560 ;
        RECT 109.685 201.390 109.855 201.580 ;
        RECT 110.150 201.390 110.320 201.580 ;
        RECT 113.360 201.390 113.530 201.580 ;
        RECT 114.745 201.390 114.915 201.580 ;
        RECT 117.515 201.415 117.675 201.525 ;
        RECT 117.960 201.420 118.080 201.530 ;
        RECT 118.425 201.370 118.595 201.560 ;
        RECT 122.105 201.370 122.275 201.560 ;
        RECT 125.335 201.415 125.495 201.525 ;
        RECT 126.250 201.370 126.420 201.560 ;
        RECT 127.165 201.390 127.335 201.580 ;
        RECT 129.465 201.560 129.615 201.580 ;
        RECT 129.465 201.390 129.635 201.560 ;
        RECT 129.935 201.415 130.095 201.525 ;
        RECT 134.065 201.370 134.235 201.560 ;
        RECT 134.525 201.370 134.695 201.560 ;
        RECT 137.285 201.370 137.455 201.560 ;
        RECT 138.670 201.370 138.840 201.560 ;
        RECT 139.125 201.390 139.295 201.580 ;
        RECT 139.585 201.390 139.755 201.580 ;
        RECT 140.965 201.530 141.135 201.560 ;
        RECT 140.055 201.415 140.215 201.525 ;
        RECT 140.960 201.420 141.135 201.530 ;
        RECT 140.965 201.370 141.135 201.420 ;
        RECT 141.425 201.390 141.595 201.580 ;
        RECT 142.805 201.390 142.975 201.580 ;
        RECT 143.265 201.370 143.435 201.560 ;
        RECT 144.645 201.370 144.815 201.580 ;
        RECT 147.405 201.370 147.575 201.580 ;
        RECT 72.700 201.340 73.655 201.370 ;
        RECT 68.835 200.460 71.225 201.140 ;
        RECT 71.375 200.660 73.655 201.340 ;
        RECT 72.700 200.460 73.655 200.660 ;
        RECT 74.585 200.460 77.795 201.370 ;
        RECT 77.805 200.460 80.725 201.370 ;
        RECT 81.655 200.460 85.155 201.370 ;
        RECT 85.165 200.460 87.775 201.370 ;
        RECT 88.380 201.140 90.070 201.370 ;
        RECT 88.380 200.460 90.215 201.140 ;
        RECT 91.155 200.500 91.585 201.285 ;
        RECT 91.685 201.140 94.675 201.370 ;
        RECT 91.685 200.460 94.745 201.140 ;
        RECT 94.825 200.560 96.655 201.370 ;
        RECT 97.125 200.460 100.335 201.370 ;
        RECT 100.345 200.560 101.715 201.370 ;
        RECT 101.725 200.460 103.075 201.370 ;
        RECT 103.105 200.460 104.455 201.370 ;
        RECT 104.485 200.460 107.695 201.370 ;
        RECT 107.705 200.690 116.810 201.370 ;
        RECT 116.915 200.500 117.345 201.285 ;
        RECT 118.395 200.690 121.860 201.370 ;
        RECT 120.940 200.460 121.860 200.690 ;
        RECT 121.965 200.460 125.175 201.370 ;
        RECT 126.105 200.690 129.690 201.370 ;
        RECT 130.800 200.690 134.265 201.370 ;
        RECT 134.385 200.690 137.135 201.370 ;
        RECT 126.105 200.460 127.025 200.690 ;
        RECT 130.800 200.460 131.720 200.690 ;
        RECT 136.205 200.460 137.135 200.690 ;
        RECT 137.155 200.460 138.505 201.370 ;
        RECT 138.525 200.460 139.875 201.370 ;
        RECT 140.825 200.690 142.655 201.370 ;
        RECT 141.310 200.460 142.655 200.690 ;
        RECT 142.675 200.500 143.105 201.285 ;
        RECT 143.135 200.460 144.485 201.370 ;
        RECT 144.505 200.690 146.335 201.370 ;
        RECT 144.990 200.460 146.335 200.690 ;
        RECT 146.345 200.560 147.715 201.370 ;
      LAYER nwell ;
        RECT 13.670 197.340 147.910 200.170 ;
      LAYER pwell ;
        RECT 13.865 196.140 15.235 196.950 ;
        RECT 15.245 196.820 16.590 197.050 ;
        RECT 22.055 196.820 22.985 197.040 ;
        RECT 25.815 196.820 26.735 197.050 ;
        RECT 15.245 196.140 17.075 196.820 ;
        RECT 17.545 196.140 26.735 196.820 ;
        RECT 26.755 196.225 27.185 197.010 ;
        RECT 27.215 196.140 29.945 197.050 ;
        RECT 29.965 196.820 31.310 197.050 ;
        RECT 29.965 196.140 31.795 196.820 ;
        RECT 32.000 196.140 35.475 197.050 ;
        RECT 35.495 196.140 38.225 197.050 ;
        RECT 38.245 196.850 39.200 197.050 ;
        RECT 38.245 196.170 40.525 196.850 ;
        RECT 38.245 196.140 39.200 196.170 ;
        RECT 14.005 195.930 14.175 196.140 ;
        RECT 16.765 195.930 16.935 196.140 ;
        RECT 17.220 195.980 17.340 196.090 ;
        RECT 17.685 195.950 17.855 196.140 ;
        RECT 18.605 195.930 18.775 196.120 ;
        RECT 19.065 195.930 19.235 196.120 ;
        RECT 27.345 195.950 27.515 196.140 ;
        RECT 31.485 195.950 31.655 196.140 ;
        RECT 32.405 195.930 32.575 196.120 ;
        RECT 13.865 195.120 15.235 195.930 ;
        RECT 15.245 195.250 17.075 195.930 ;
        RECT 17.085 195.250 18.915 195.930 ;
        RECT 18.925 195.250 29.295 195.930 ;
        RECT 15.245 195.020 16.590 195.250 ;
        RECT 17.085 195.020 18.430 195.250 ;
        RECT 23.435 195.030 24.365 195.250 ;
        RECT 27.085 195.020 29.295 195.250 ;
        RECT 29.505 195.020 32.715 195.930 ;
        RECT 32.865 195.900 33.035 196.120 ;
        RECT 35.160 195.950 35.330 196.140 ;
        RECT 35.625 195.950 35.795 196.140 ;
        RECT 36.080 195.980 36.200 196.090 ;
        RECT 36.545 195.930 36.715 196.120 ;
        RECT 39.300 195.930 39.470 196.120 ;
        RECT 40.230 195.930 40.400 196.170 ;
        RECT 41.485 196.140 42.835 197.050 ;
        RECT 43.775 196.140 46.975 197.050 ;
        RECT 46.995 196.140 50.195 197.050 ;
        RECT 50.205 196.140 51.555 197.050 ;
        RECT 52.515 196.225 52.945 197.010 ;
        RECT 52.965 196.140 54.335 196.920 ;
        RECT 54.345 196.140 55.715 196.950 ;
        RECT 55.735 196.140 57.085 197.050 ;
        RECT 57.125 196.140 58.475 197.050 ;
        RECT 58.485 196.140 59.835 197.050 ;
        RECT 64.375 196.820 65.305 197.040 ;
        RECT 68.025 196.820 70.235 197.050 ;
        RECT 72.520 196.820 73.655 197.050 ;
        RECT 75.035 196.820 75.955 197.050 ;
        RECT 59.865 196.140 70.235 196.820 ;
        RECT 70.445 196.140 73.655 196.820 ;
        RECT 73.665 196.140 75.955 196.820 ;
        RECT 76.425 196.820 77.770 197.050 ;
        RECT 76.425 196.140 78.255 196.820 ;
        RECT 78.275 196.225 78.705 197.010 ;
        RECT 78.725 196.140 81.935 197.050 ;
        RECT 83.045 196.370 85.380 197.050 ;
        RECT 83.045 196.140 84.895 196.370 ;
        RECT 85.625 196.140 89.295 196.950 ;
        RECT 89.305 196.140 90.675 196.950 ;
        RECT 90.705 196.140 92.055 197.050 ;
        RECT 92.065 196.140 97.575 196.950 ;
        RECT 100.120 196.820 101.255 197.050 ;
        RECT 98.045 196.140 101.255 196.820 ;
        RECT 101.500 196.370 103.835 197.050 ;
        RECT 101.985 196.140 103.835 196.370 ;
        RECT 104.035 196.225 104.465 197.010 ;
        RECT 106.560 196.820 107.695 197.050 ;
        RECT 104.485 196.140 107.695 196.820 ;
        RECT 107.705 196.850 108.635 197.050 ;
        RECT 109.965 196.850 110.915 197.050 ;
        RECT 107.705 196.370 110.915 196.850 ;
        RECT 115.435 196.820 116.365 197.040 ;
        RECT 119.085 196.820 121.295 197.050 ;
        RECT 107.850 196.170 110.915 196.370 ;
        RECT 40.695 195.985 40.855 196.095 ;
        RECT 41.600 195.950 41.770 196.140 ;
        RECT 42.995 195.985 43.155 196.095 ;
        RECT 43.900 195.950 44.070 196.140 ;
        RECT 34.990 195.900 35.935 195.930 ;
        RECT 32.865 195.700 35.935 195.900 ;
        RECT 32.725 195.220 35.935 195.700 ;
        RECT 32.725 195.020 33.655 195.220 ;
        RECT 34.990 195.020 35.935 195.220 ;
        RECT 36.415 195.020 37.765 195.930 ;
        RECT 37.845 195.020 39.615 195.930 ;
        RECT 39.635 195.060 40.065 195.845 ;
        RECT 40.085 195.020 43.955 195.930 ;
        RECT 44.360 195.900 44.530 196.120 ;
        RECT 47.120 195.950 47.290 196.140 ;
        RECT 47.590 195.930 47.760 196.120 ;
        RECT 51.270 195.950 51.440 196.140 ;
        RECT 51.450 195.930 51.620 196.120 ;
        RECT 51.735 195.985 51.895 196.095 ;
        RECT 52.190 195.930 52.360 196.120 ;
        RECT 54.025 195.950 54.195 196.140 ;
        RECT 54.485 195.950 54.655 196.140 ;
        RECT 55.405 195.930 55.575 196.120 ;
        RECT 56.785 195.950 56.955 196.140 ;
        RECT 57.240 195.950 57.410 196.140 ;
        RECT 58.625 195.930 58.795 196.120 ;
        RECT 59.550 195.950 59.720 196.140 ;
        RECT 60.005 195.950 60.175 196.140 ;
        RECT 61.845 195.930 62.015 196.120 ;
        RECT 65.985 195.930 66.155 196.120 ;
        RECT 69.205 195.930 69.375 196.120 ;
        RECT 70.585 195.950 70.755 196.140 ;
        RECT 73.805 195.950 73.975 196.140 ;
        RECT 76.100 195.980 76.220 196.090 ;
        RECT 77.945 195.950 78.115 196.140 ;
        RECT 78.865 195.950 79.035 196.140 ;
        RECT 83.045 196.120 83.175 196.140 ;
        RECT 82.095 195.985 82.255 196.095 ;
        RECT 83.005 195.950 83.175 196.120 ;
        RECT 85.765 195.950 85.935 196.140 ;
        RECT 89.445 195.950 89.615 196.140 ;
        RECT 91.740 196.120 91.910 196.140 ;
        RECT 89.905 195.930 90.075 196.120 ;
        RECT 90.375 195.975 90.535 196.085 ;
        RECT 91.740 195.950 91.915 196.120 ;
        RECT 92.205 195.950 92.375 196.140 ;
        RECT 97.720 195.980 97.840 196.090 ;
        RECT 98.185 195.950 98.355 196.140 ;
        RECT 103.705 196.120 103.835 196.140 ;
        RECT 91.745 195.930 91.915 195.950 ;
        RECT 103.245 195.930 103.415 196.120 ;
        RECT 103.705 195.950 103.880 196.120 ;
        RECT 104.625 195.950 104.795 196.140 ;
        RECT 105.095 195.975 105.255 196.085 ;
        RECT 103.710 195.930 103.880 195.950 ;
        RECT 106.925 195.930 107.095 196.120 ;
        RECT 107.850 195.950 108.020 196.170 ;
        RECT 109.980 196.140 110.915 196.170 ;
        RECT 110.925 196.140 121.295 196.820 ;
        RECT 121.600 196.820 122.520 197.050 ;
        RECT 121.600 196.140 125.065 196.820 ;
        RECT 125.185 196.140 127.935 197.050 ;
        RECT 127.945 196.820 129.290 197.050 ;
        RECT 127.945 196.140 129.775 196.820 ;
        RECT 129.795 196.225 130.225 197.010 ;
        RECT 131.215 196.140 135.685 197.050 ;
        RECT 135.765 196.140 137.135 196.920 ;
        RECT 137.630 196.820 138.975 197.050 ;
        RECT 139.470 196.820 140.815 197.050 ;
        RECT 141.310 196.820 142.655 197.050 ;
        RECT 143.150 196.820 144.495 197.050 ;
        RECT 144.990 196.820 146.335 197.050 ;
        RECT 137.145 196.140 138.975 196.820 ;
        RECT 138.985 196.140 140.815 196.820 ;
        RECT 140.825 196.140 142.655 196.820 ;
        RECT 142.665 196.140 144.495 196.820 ;
        RECT 144.505 196.140 146.335 196.820 ;
        RECT 146.345 196.140 147.715 196.950 ;
        RECT 110.145 195.930 110.315 196.120 ;
        RECT 110.600 195.980 110.720 196.090 ;
        RECT 111.065 195.950 111.235 196.140 ;
        RECT 113.365 195.930 113.535 196.120 ;
        RECT 113.825 195.930 113.995 196.120 ;
        RECT 117.505 195.950 117.675 196.120 ;
        RECT 117.545 195.930 117.675 195.950 ;
        RECT 120.265 195.930 120.435 196.120 ;
        RECT 124.865 195.950 125.035 196.140 ;
        RECT 127.625 195.950 127.795 196.140 ;
        RECT 129.465 196.120 129.635 196.140 ;
        RECT 129.465 195.950 129.640 196.120 ;
        RECT 130.395 195.985 130.555 196.095 ;
        RECT 131.285 195.950 131.455 196.140 ;
        RECT 129.470 195.930 129.640 195.950 ;
        RECT 135.905 195.930 136.075 196.120 ;
        RECT 136.825 195.950 136.995 196.140 ;
        RECT 137.285 195.950 137.455 196.140 ;
        RECT 137.745 195.930 137.915 196.120 ;
        RECT 138.205 195.930 138.375 196.120 ;
        RECT 139.125 195.950 139.295 196.140 ;
        RECT 140.055 195.975 140.215 196.085 ;
        RECT 140.965 195.930 141.135 196.140 ;
        RECT 142.805 195.950 142.975 196.140 ;
        RECT 143.270 195.930 143.440 196.120 ;
        RECT 144.645 195.930 144.815 196.140 ;
        RECT 147.405 195.930 147.575 196.140 ;
        RECT 45.560 195.900 46.515 195.930 ;
        RECT 44.235 195.220 46.515 195.900 ;
        RECT 45.560 195.020 46.515 195.220 ;
        RECT 46.525 195.020 47.875 195.930 ;
        RECT 48.135 195.250 52.035 195.930 ;
        RECT 51.105 195.020 52.035 195.250 ;
        RECT 52.045 195.020 54.965 195.930 ;
        RECT 55.265 195.020 58.475 195.930 ;
        RECT 58.485 195.020 61.695 195.930 ;
        RECT 61.705 195.120 65.375 195.930 ;
        RECT 65.395 195.060 65.825 195.845 ;
        RECT 65.845 195.020 69.055 195.930 ;
        RECT 69.065 195.250 79.435 195.930 ;
        RECT 73.575 195.030 74.505 195.250 ;
        RECT 77.225 195.020 79.435 195.250 ;
        RECT 79.845 195.250 90.215 195.930 ;
        RECT 79.845 195.020 82.055 195.250 ;
        RECT 84.775 195.030 85.705 195.250 ;
        RECT 91.155 195.060 91.585 195.845 ;
        RECT 91.605 195.250 101.975 195.930 ;
        RECT 96.115 195.030 97.045 195.250 ;
        RECT 99.765 195.020 101.975 195.250 ;
        RECT 102.185 195.150 103.555 195.930 ;
        RECT 103.565 195.020 104.915 195.930 ;
        RECT 105.865 195.150 107.235 195.930 ;
        RECT 107.245 195.020 110.415 195.930 ;
        RECT 110.935 195.020 113.665 195.930 ;
        RECT 113.685 195.020 116.895 195.930 ;
        RECT 116.915 195.060 117.345 195.845 ;
        RECT 117.545 195.700 119.395 195.930 ;
        RECT 117.545 195.020 119.880 195.700 ;
        RECT 120.125 195.250 129.315 195.930 ;
        RECT 124.635 195.030 125.565 195.250 ;
        RECT 128.395 195.020 129.315 195.250 ;
        RECT 129.325 195.020 133.455 195.930 ;
        RECT 133.475 195.020 136.205 195.930 ;
        RECT 136.225 195.250 138.055 195.930 ;
        RECT 138.065 195.250 139.895 195.930 ;
        RECT 140.825 195.250 142.655 195.930 ;
        RECT 136.225 195.020 137.570 195.250 ;
        RECT 138.550 195.020 139.895 195.250 ;
        RECT 141.310 195.020 142.655 195.250 ;
        RECT 142.675 195.060 143.105 195.845 ;
        RECT 143.125 195.020 144.475 195.930 ;
        RECT 144.505 195.250 146.335 195.930 ;
        RECT 144.990 195.020 146.335 195.250 ;
        RECT 146.345 195.120 147.715 195.930 ;
      LAYER nwell ;
        RECT 13.670 191.900 147.910 194.730 ;
      LAYER pwell ;
        RECT 13.865 190.700 15.235 191.510 ;
        RECT 15.245 191.380 16.590 191.610 ;
        RECT 17.085 191.380 18.430 191.610 ;
        RECT 18.925 191.380 20.270 191.610 ;
        RECT 20.765 191.380 22.110 191.610 ;
        RECT 25.390 191.380 26.735 191.610 ;
        RECT 15.245 190.700 17.075 191.380 ;
        RECT 17.085 190.700 18.915 191.380 ;
        RECT 18.925 190.700 20.755 191.380 ;
        RECT 20.765 190.700 22.595 191.380 ;
        RECT 23.065 190.700 24.895 191.380 ;
        RECT 24.905 190.700 26.735 191.380 ;
        RECT 26.755 190.785 27.185 191.570 ;
        RECT 27.205 190.700 30.415 191.610 ;
        RECT 30.425 191.380 31.770 191.610 ;
        RECT 32.265 191.380 33.610 191.610 ;
        RECT 34.105 191.410 35.035 191.610 ;
        RECT 36.370 191.410 37.315 191.610 ;
        RECT 30.425 190.700 32.255 191.380 ;
        RECT 32.265 190.700 34.095 191.380 ;
        RECT 34.105 190.930 37.315 191.410 ;
        RECT 34.245 190.730 37.315 190.930 ;
        RECT 14.005 190.510 14.175 190.700 ;
        RECT 16.765 190.510 16.935 190.700 ;
        RECT 18.605 190.510 18.775 190.700 ;
        RECT 20.445 190.510 20.615 190.700 ;
        RECT 22.285 190.510 22.455 190.700 ;
        RECT 22.740 190.540 22.860 190.650 ;
        RECT 23.205 190.510 23.375 190.700 ;
        RECT 25.045 190.510 25.215 190.700 ;
        RECT 30.105 190.510 30.275 190.700 ;
        RECT 31.945 190.510 32.115 190.700 ;
        RECT 33.785 190.510 33.955 190.700 ;
        RECT 34.245 190.510 34.415 190.730 ;
        RECT 36.370 190.700 37.315 190.730 ;
        RECT 37.325 191.380 38.670 191.610 ;
        RECT 37.325 190.700 39.155 191.380 ;
        RECT 39.635 190.785 40.065 191.570 ;
        RECT 40.085 190.700 41.455 191.480 ;
        RECT 41.465 190.700 42.835 191.480 ;
        RECT 42.865 190.700 44.215 191.610 ;
        RECT 44.710 191.380 46.055 191.610 ;
        RECT 44.225 190.700 46.055 191.380 ;
        RECT 46.300 190.930 48.635 191.610 ;
        RECT 46.785 190.700 48.635 190.930 ;
        RECT 48.825 190.700 52.035 191.610 ;
        RECT 52.515 190.785 52.945 191.570 ;
        RECT 53.905 190.700 55.255 191.610 ;
        RECT 55.905 190.930 58.240 191.610 ;
        RECT 58.970 191.380 60.315 191.610 ;
        RECT 55.905 190.700 57.755 190.930 ;
        RECT 58.485 190.700 60.315 191.380 ;
        RECT 60.325 190.700 61.695 191.480 ;
        RECT 61.705 190.700 63.055 191.610 ;
        RECT 63.105 190.700 64.455 191.610 ;
        RECT 65.395 190.785 65.825 191.570 ;
        RECT 66.330 191.380 67.675 191.610 ;
        RECT 65.845 190.700 67.675 191.380 ;
        RECT 67.685 190.700 69.515 191.510 ;
        RECT 69.525 190.700 70.895 191.480 ;
        RECT 70.925 190.700 72.275 191.610 ;
        RECT 72.285 190.700 73.655 191.480 ;
        RECT 74.150 191.380 75.495 191.610 ;
        RECT 73.665 190.700 75.495 191.380 ;
        RECT 75.685 190.930 78.020 191.610 ;
        RECT 75.685 190.700 77.535 190.930 ;
        RECT 78.275 190.785 78.705 191.570 ;
        RECT 78.725 190.700 81.935 191.610 ;
        RECT 81.965 190.700 83.315 191.610 ;
        RECT 83.810 191.380 85.155 191.610 ;
        RECT 83.325 190.700 85.155 191.380 ;
        RECT 86.085 190.700 87.455 191.480 ;
        RECT 87.465 190.700 90.675 191.610 ;
        RECT 91.155 190.785 91.585 191.570 ;
        RECT 93.010 191.380 94.355 191.610 ;
        RECT 92.525 190.700 94.355 191.380 ;
        RECT 95.060 190.930 97.395 191.610 ;
        RECT 95.545 190.700 97.395 190.930 ;
        RECT 97.585 190.700 100.795 191.610 ;
        RECT 101.725 191.380 103.070 191.610 ;
        RECT 101.725 190.700 103.555 191.380 ;
        RECT 104.035 190.785 104.465 191.570 ;
        RECT 104.685 191.380 106.895 191.610 ;
        RECT 109.615 191.380 110.545 191.600 ;
        RECT 115.065 191.380 116.410 191.610 ;
        RECT 104.685 190.700 115.055 191.380 ;
        RECT 115.065 190.700 116.895 191.380 ;
        RECT 116.915 190.785 117.345 191.570 ;
        RECT 117.365 190.700 118.735 191.480 ;
        RECT 119.665 190.700 123.335 191.610 ;
        RECT 125.165 191.380 126.095 191.610 ;
        RECT 123.345 190.700 126.095 191.380 ;
        RECT 126.105 191.380 127.450 191.610 ;
        RECT 128.430 191.380 129.775 191.610 ;
        RECT 126.105 190.700 127.935 191.380 ;
        RECT 127.945 190.700 129.775 191.380 ;
        RECT 129.795 190.785 130.225 191.570 ;
        RECT 130.730 191.380 132.075 191.610 ;
        RECT 130.245 190.700 132.075 191.380 ;
        RECT 133.005 191.380 134.350 191.610 ;
        RECT 133.005 190.700 134.835 191.380 ;
        RECT 134.865 190.700 136.215 191.610 ;
        RECT 137.365 191.520 138.315 191.610 ;
        RECT 140.125 191.520 141.075 191.610 ;
        RECT 136.385 190.700 138.315 191.520 ;
        RECT 139.145 190.700 141.075 191.520 ;
        RECT 141.285 190.700 142.635 191.610 ;
        RECT 142.675 190.785 143.105 191.570 ;
        RECT 143.585 190.700 146.325 191.380 ;
        RECT 146.345 190.700 147.715 191.510 ;
        RECT 38.845 190.510 39.015 190.700 ;
        RECT 39.300 190.540 39.420 190.650 ;
        RECT 41.145 190.510 41.315 190.700 ;
        RECT 41.605 190.510 41.775 190.700 ;
        RECT 43.900 190.510 44.070 190.700 ;
        RECT 44.365 190.510 44.535 190.700 ;
        RECT 48.505 190.680 48.635 190.700 ;
        RECT 48.505 190.510 48.675 190.680 ;
        RECT 48.965 190.510 49.135 190.700 ;
        RECT 52.180 190.540 52.300 190.650 ;
        RECT 53.115 190.545 53.275 190.655 ;
        RECT 54.940 190.510 55.110 190.700 ;
        RECT 55.905 190.680 56.035 190.700 ;
        RECT 55.400 190.540 55.520 190.650 ;
        RECT 55.865 190.510 56.035 190.680 ;
        RECT 58.625 190.510 58.795 190.700 ;
        RECT 61.385 190.510 61.555 190.700 ;
        RECT 61.850 190.510 62.020 190.700 ;
        RECT 64.140 190.510 64.310 190.700 ;
        RECT 64.615 190.545 64.775 190.655 ;
        RECT 65.985 190.510 66.155 190.700 ;
        RECT 67.825 190.510 67.995 190.700 ;
        RECT 69.665 190.510 69.835 190.700 ;
        RECT 71.960 190.510 72.130 190.700 ;
        RECT 72.425 190.510 72.595 190.700 ;
        RECT 73.805 190.510 73.975 190.700 ;
        RECT 75.685 190.680 75.815 190.700 ;
        RECT 75.645 190.510 75.815 190.680 ;
        RECT 78.865 190.510 79.035 190.700 ;
        RECT 83.000 190.510 83.170 190.700 ;
        RECT 83.465 190.510 83.635 190.700 ;
        RECT 85.315 190.545 85.475 190.655 ;
        RECT 87.145 190.510 87.315 190.700 ;
        RECT 87.605 190.510 87.775 190.700 ;
        RECT 90.820 190.540 90.940 190.650 ;
        RECT 91.755 190.545 91.915 190.655 ;
        RECT 92.665 190.510 92.835 190.700 ;
        RECT 97.265 190.680 97.395 190.700 ;
        RECT 94.500 190.540 94.620 190.650 ;
        RECT 97.265 190.510 97.435 190.680 ;
        RECT 97.725 190.510 97.895 190.700 ;
        RECT 100.955 190.545 101.115 190.655 ;
        RECT 103.245 190.510 103.415 190.700 ;
        RECT 103.700 190.540 103.820 190.650 ;
        RECT 114.745 190.510 114.915 190.700 ;
        RECT 116.585 190.510 116.755 190.700 ;
        RECT 117.505 190.510 117.675 190.700 ;
        RECT 118.895 190.545 119.055 190.655 ;
        RECT 119.810 190.510 119.980 190.700 ;
        RECT 123.485 190.510 123.655 190.700 ;
        RECT 127.625 190.510 127.795 190.700 ;
        RECT 128.085 190.510 128.255 190.700 ;
        RECT 130.385 190.510 130.555 190.700 ;
        RECT 132.235 190.545 132.395 190.655 ;
        RECT 134.525 190.510 134.695 190.700 ;
        RECT 135.900 190.510 136.070 190.700 ;
        RECT 136.385 190.680 136.535 190.700 ;
        RECT 139.145 190.680 139.295 190.700 ;
        RECT 136.365 190.510 136.535 190.680 ;
        RECT 138.660 190.540 138.780 190.650 ;
        RECT 139.125 190.510 139.295 190.680 ;
        RECT 141.430 190.510 141.600 190.700 ;
        RECT 143.260 190.540 143.380 190.650 ;
        RECT 143.725 190.510 143.895 190.700 ;
        RECT 147.405 190.510 147.575 190.700 ;
      LAYER nwell ;
        RECT 109.245 183.595 141.785 185.365 ;
      LAYER pwell ;
        RECT 142.880 184.815 143.050 184.985 ;
        RECT 142.880 184.795 142.985 184.815 ;
        RECT 144.265 184.795 144.435 184.985 ;
        RECT 142.055 183.885 142.985 184.795 ;
        RECT 143.200 183.885 144.550 184.795 ;
        RECT 8.180 182.470 8.350 182.660 ;
        RECT 11.400 182.470 11.570 182.660 ;
        RECT 16.920 182.470 17.090 182.660 ;
        RECT 18.305 182.470 18.475 182.660 ;
        RECT 8.040 181.560 11.225 182.470 ;
        RECT 11.260 181.660 16.770 182.470 ;
        RECT 16.780 181.660 18.150 182.470 ;
        RECT 18.160 181.560 21.275 182.470 ;
      LAYER nwell ;
        RECT 7.845 178.440 21.565 181.270 ;
        RECT 39.270 180.030 46.120 180.070 ;
        RECT 35.400 178.425 46.120 180.030 ;
      LAYER pwell ;
        RECT 8.040 177.240 11.225 178.150 ;
        RECT 11.260 177.240 14.445 178.150 ;
        RECT 14.490 177.325 14.920 178.110 ;
        RECT 14.940 177.240 18.055 178.150 ;
        RECT 18.160 177.240 21.275 178.150 ;
        RECT 8.180 177.030 8.350 177.240 ;
        RECT 11.400 177.030 11.570 177.240 ;
        RECT 15.085 177.030 15.255 177.240 ;
        RECT 18.305 177.030 18.475 177.240 ;
        RECT 35.645 177.225 37.835 178.135 ;
        RECT 38.130 177.225 39.060 178.135 ;
        RECT 8.040 176.120 11.225 177.030 ;
        RECT 11.260 176.120 14.445 177.030 ;
        RECT 14.490 176.160 14.920 176.945 ;
        RECT 14.940 176.120 18.055 177.030 ;
        RECT 18.160 176.120 21.275 177.030 ;
        RECT 37.575 177.015 37.745 177.225 ;
        RECT 38.955 177.205 39.060 177.225 ;
        RECT 38.955 177.035 39.125 177.205 ;
        RECT 38.955 177.015 39.060 177.035 ;
        RECT 35.645 176.105 37.835 177.015 ;
        RECT 38.130 176.105 39.060 177.015 ;
      LAYER nwell ;
        RECT 7.845 173.000 21.565 175.830 ;
        RECT 39.270 175.815 46.120 178.425 ;
        RECT 35.400 173.880 46.120 175.815 ;
      LAYER pwell ;
        RECT 47.780 178.100 71.600 181.120 ;
      LAYER nwell ;
        RECT 71.600 181.110 73.710 181.120 ;
        RECT 71.600 178.280 102.600 181.110 ;
        RECT 35.400 172.985 38.540 173.880 ;
      LAYER pwell ;
        RECT 8.040 171.800 11.225 172.710 ;
        RECT 11.260 171.800 14.445 172.710 ;
        RECT 14.490 171.885 14.920 172.670 ;
        RECT 14.940 171.800 18.055 172.710 ;
        RECT 18.160 171.800 21.275 172.710 ;
        RECT 8.180 171.590 8.350 171.800 ;
        RECT 11.400 171.590 11.570 171.800 ;
        RECT 15.085 171.590 15.255 171.800 ;
        RECT 18.305 171.590 18.475 171.800 ;
        RECT 35.595 171.785 38.205 172.695 ;
        RECT 35.740 171.595 35.910 171.785 ;
        RECT 8.040 170.680 11.225 171.590 ;
        RECT 11.260 170.680 14.445 171.590 ;
        RECT 14.490 170.720 14.920 171.505 ;
        RECT 14.940 170.680 18.055 171.590 ;
        RECT 18.160 170.680 21.275 171.590 ;
        RECT 39.275 170.780 46.125 173.880 ;
        RECT 47.780 170.810 73.710 178.100 ;
      LAYER nwell ;
        RECT 73.710 170.960 102.600 178.280 ;
        RECT 109.245 180.765 144.765 183.595 ;
        RECT 109.245 178.155 141.785 180.765 ;
      LAYER pwell ;
        RECT 142.055 179.565 142.985 180.475 ;
        RECT 143.200 179.565 144.550 180.475 ;
        RECT 142.880 179.545 142.985 179.565 ;
        RECT 142.880 179.375 143.050 179.545 ;
        RECT 144.265 179.375 144.435 179.565 ;
        RECT 142.880 179.355 142.985 179.375 ;
        RECT 144.715 179.355 144.885 179.545 ;
        RECT 142.055 178.445 142.985 179.355 ;
        RECT 143.200 178.445 145.030 179.355 ;
      LAYER nwell ;
        RECT 109.245 176.550 145.225 178.155 ;
        RECT 109.245 175.325 144.765 176.550 ;
        RECT 109.245 172.835 141.785 175.325 ;
      LAYER pwell ;
        RECT 142.025 174.125 142.955 175.035 ;
        RECT 143.405 174.125 144.335 175.035 ;
        RECT 142.025 174.105 142.130 174.125 ;
        RECT 143.405 174.105 143.510 174.125 ;
        RECT 141.960 173.935 142.130 174.105 ;
        RECT 143.340 173.935 143.510 174.105 ;
      LAYER nwell ;
        RECT 73.710 170.920 102.610 170.960 ;
        RECT 7.845 167.560 21.565 170.390 ;
      LAYER pwell ;
        RECT 39.275 170.310 41.385 170.780 ;
        RECT 44.015 170.310 46.125 170.780 ;
        RECT 39.275 169.780 46.125 170.310 ;
        RECT 8.040 166.360 11.225 167.270 ;
        RECT 11.260 166.360 14.445 167.270 ;
        RECT 14.490 166.445 14.920 167.230 ;
        RECT 14.940 166.360 18.055 167.270 ;
        RECT 18.160 166.360 21.275 167.270 ;
        RECT 40.010 167.210 45.310 169.780 ;
        RECT 8.180 166.170 8.350 166.360 ;
        RECT 11.400 166.170 11.570 166.360 ;
        RECT 15.085 166.170 15.255 166.360 ;
        RECT 18.305 166.170 18.475 166.360 ;
        RECT 47.780 165.740 54.430 169.840 ;
      LAYER nwell ;
        RECT 54.590 165.740 61.240 169.930 ;
      LAYER pwell ;
        RECT 62.880 165.740 66.470 169.740 ;
        RECT 71.600 168.510 73.710 170.810 ;
        RECT 68.090 165.740 73.710 168.510 ;
      LAYER nwell ;
        RECT 73.710 165.740 84.360 170.920 ;
      LAYER pwell ;
        RECT 84.490 166.700 90.840 170.800 ;
      LAYER nwell ;
        RECT 91.730 168.610 95.980 170.920 ;
        RECT 100.850 169.355 102.610 170.920 ;
      LAYER pwell ;
        RECT 101.280 168.155 102.210 169.065 ;
        RECT 102.105 168.135 102.210 168.155 ;
      LAYER nwell ;
        RECT 109.245 168.145 144.845 172.835 ;
      LAYER pwell ;
        RECT 102.105 167.965 102.275 168.135 ;
      LAYER nwell ;
        RECT 109.245 161.515 141.785 168.145 ;
      LAYER pwell ;
        RECT 141.795 162.675 144.905 167.185 ;
        RECT 20.260 160.210 24.000 160.215 ;
        RECT 30.815 160.210 37.715 160.270 ;
        RECT 123.400 160.210 130.300 160.270 ;
        RECT 137.115 160.210 140.855 160.215 ;
        RECT 20.260 159.955 37.715 160.210 ;
        RECT 22.190 159.840 22.360 159.955 ;
        RECT 22.425 159.840 37.715 159.955 ;
        RECT 20.260 158.930 37.715 159.840 ;
      LAYER nwell ;
        RECT 20.015 156.280 24.075 158.640 ;
        RECT 20.010 155.810 24.075 156.280 ;
        RECT 20.010 155.095 21.335 155.810 ;
      LAYER pwell ;
        RECT 24.075 155.520 37.715 158.930 ;
        RECT 21.640 154.110 37.715 155.520 ;
        RECT 30.815 153.690 37.715 154.110 ;
      LAYER nwell ;
        RECT 37.715 154.020 74.605 160.210 ;
        RECT 40.720 154.015 74.605 154.020 ;
        RECT 42.275 149.365 74.605 154.015 ;
        RECT 42.355 149.340 74.605 149.365 ;
        RECT 86.510 154.020 123.400 160.210 ;
      LAYER pwell ;
        RECT 123.400 159.955 140.855 160.210 ;
        RECT 123.400 159.840 138.690 159.955 ;
        RECT 138.755 159.840 138.925 159.955 ;
        RECT 123.400 158.930 140.855 159.840 ;
        RECT 123.400 155.520 137.040 158.930 ;
      LAYER nwell ;
        RECT 137.040 156.280 141.100 158.640 ;
        RECT 137.040 155.810 141.105 156.280 ;
      LAYER pwell ;
        RECT 123.400 154.110 139.475 155.520 ;
      LAYER nwell ;
        RECT 139.780 155.095 141.105 155.810 ;
        RECT 86.510 154.015 120.395 154.020 ;
        RECT 86.510 149.365 118.840 154.015 ;
      LAYER pwell ;
        RECT 123.400 153.690 130.300 154.110 ;
      LAYER nwell ;
        RECT 86.510 149.340 118.760 149.365 ;
        RECT 7.285 133.075 36.095 142.915 ;
      LAYER pwell ;
        RECT 36.105 133.075 75.325 142.925 ;
        RECT 85.790 133.075 125.010 142.925 ;
      LAYER nwell ;
        RECT 125.020 133.075 153.830 142.915 ;
      LAYER pwell ;
        RECT 6.840 4.990 74.540 126.640 ;
        RECT 86.575 4.990 154.275 126.640 ;
      LAYER li1 ;
        RECT 13.860 217.710 147.720 217.880 ;
        RECT 13.945 216.960 15.155 217.710 ;
        RECT 15.385 217.230 15.665 217.710 ;
        RECT 15.835 217.060 16.095 217.450 ;
        RECT 16.270 217.230 16.525 217.710 ;
        RECT 16.695 217.060 16.990 217.450 ;
        RECT 17.170 217.230 17.445 217.710 ;
        RECT 17.615 217.210 17.915 217.540 ;
        RECT 13.945 216.420 14.465 216.960 ;
        RECT 15.340 216.890 16.990 217.060 ;
        RECT 14.635 216.250 15.155 216.790 ;
        RECT 13.945 215.160 15.155 216.250 ;
        RECT 15.340 216.380 15.745 216.890 ;
        RECT 15.915 216.550 17.055 216.720 ;
        RECT 15.340 216.210 16.095 216.380 ;
        RECT 15.380 215.160 15.665 216.030 ;
        RECT 15.835 215.960 16.095 216.210 ;
        RECT 16.885 216.300 17.055 216.550 ;
        RECT 17.225 216.470 17.575 217.040 ;
        RECT 17.745 216.300 17.915 217.210 ;
        RECT 18.090 216.870 18.350 217.710 ;
        RECT 18.525 216.965 18.780 217.540 ;
        RECT 18.950 217.330 19.280 217.710 ;
        RECT 19.495 217.160 19.665 217.540 ;
        RECT 18.950 216.990 19.665 217.160 ;
        RECT 16.885 216.130 17.915 216.300 ;
        RECT 15.835 215.790 16.955 215.960 ;
        RECT 15.835 215.330 16.095 215.790 ;
        RECT 16.270 215.160 16.525 215.620 ;
        RECT 16.695 215.330 16.955 215.790 ;
        RECT 17.125 215.160 17.435 215.960 ;
        RECT 17.605 215.330 17.915 216.130 ;
        RECT 18.090 215.160 18.350 216.310 ;
        RECT 18.525 216.235 18.695 216.965 ;
        RECT 18.950 216.800 19.120 216.990 ;
        RECT 19.930 216.870 20.190 217.710 ;
        RECT 20.365 216.965 20.620 217.540 ;
        RECT 20.790 217.330 21.120 217.710 ;
        RECT 21.335 217.160 21.505 217.540 ;
        RECT 20.790 216.990 21.505 217.160 ;
        RECT 21.855 217.160 22.025 217.540 ;
        RECT 22.205 217.330 22.535 217.710 ;
        RECT 21.855 216.990 22.520 217.160 ;
        RECT 22.715 217.035 22.975 217.540 ;
        RECT 18.865 216.470 19.120 216.800 ;
        RECT 18.950 216.260 19.120 216.470 ;
        RECT 19.400 216.440 19.755 216.810 ;
        RECT 18.525 215.330 18.780 216.235 ;
        RECT 18.950 216.090 19.665 216.260 ;
        RECT 18.950 215.160 19.280 215.920 ;
        RECT 19.495 215.330 19.665 216.090 ;
        RECT 19.930 215.160 20.190 216.310 ;
        RECT 20.365 216.235 20.535 216.965 ;
        RECT 20.790 216.800 20.960 216.990 ;
        RECT 20.705 216.470 20.960 216.800 ;
        RECT 20.790 216.260 20.960 216.470 ;
        RECT 21.240 216.440 21.595 216.810 ;
        RECT 21.785 216.440 22.125 216.810 ;
        RECT 22.350 216.735 22.520 216.990 ;
        RECT 22.350 216.405 22.625 216.735 ;
        RECT 22.350 216.260 22.520 216.405 ;
        RECT 20.365 215.330 20.620 216.235 ;
        RECT 20.790 216.090 21.505 216.260 ;
        RECT 20.790 215.160 21.120 215.920 ;
        RECT 21.335 215.330 21.505 216.090 ;
        RECT 21.845 216.090 22.520 216.260 ;
        RECT 22.795 216.235 22.975 217.035 ;
        RECT 23.145 216.940 24.815 217.710 ;
        RECT 23.145 216.420 23.895 216.940 ;
        RECT 25.505 216.890 25.715 217.710 ;
        RECT 25.885 216.910 26.215 217.540 ;
        RECT 24.065 216.250 24.815 216.770 ;
        RECT 25.885 216.310 26.135 216.910 ;
        RECT 26.385 216.890 26.615 217.710 ;
        RECT 26.825 216.985 27.115 217.710 ;
        RECT 27.290 216.970 27.545 217.540 ;
        RECT 27.715 217.310 28.045 217.710 ;
        RECT 28.470 217.175 29.000 217.540 ;
        RECT 29.190 217.370 29.465 217.540 ;
        RECT 29.185 217.200 29.465 217.370 ;
        RECT 28.470 217.140 28.645 217.175 ;
        RECT 27.715 216.970 28.645 217.140 ;
        RECT 26.305 216.470 26.635 216.720 ;
        RECT 21.845 215.330 22.025 216.090 ;
        RECT 22.205 215.160 22.535 215.920 ;
        RECT 22.705 215.330 22.975 216.235 ;
        RECT 23.145 215.160 24.815 216.250 ;
        RECT 25.505 215.160 25.715 216.300 ;
        RECT 25.885 215.330 26.215 216.310 ;
        RECT 26.385 215.160 26.615 216.300 ;
        RECT 26.825 215.160 27.115 216.325 ;
        RECT 27.290 216.300 27.460 216.970 ;
        RECT 27.715 216.800 27.885 216.970 ;
        RECT 27.630 216.470 27.885 216.800 ;
        RECT 28.110 216.470 28.305 216.800 ;
        RECT 27.290 215.330 27.625 216.300 ;
        RECT 27.795 215.160 27.965 216.300 ;
        RECT 28.135 215.500 28.305 216.470 ;
        RECT 28.475 215.840 28.645 216.970 ;
        RECT 28.815 216.180 28.985 216.980 ;
        RECT 29.190 216.380 29.465 217.200 ;
        RECT 29.635 216.180 29.825 217.540 ;
        RECT 30.005 217.175 30.515 217.710 ;
        RECT 30.735 216.900 30.980 217.505 ;
        RECT 31.425 217.210 31.725 217.540 ;
        RECT 31.895 217.230 32.170 217.710 ;
        RECT 30.025 216.730 31.255 216.900 ;
        RECT 28.815 216.010 29.825 216.180 ;
        RECT 29.995 216.165 30.745 216.355 ;
        RECT 28.475 215.670 29.600 215.840 ;
        RECT 29.995 215.500 30.165 216.165 ;
        RECT 30.915 215.920 31.255 216.730 ;
        RECT 28.135 215.330 30.165 215.500 ;
        RECT 30.335 215.160 30.505 215.920 ;
        RECT 30.740 215.510 31.255 215.920 ;
        RECT 31.425 216.300 31.595 217.210 ;
        RECT 32.350 217.060 32.645 217.450 ;
        RECT 32.815 217.230 33.070 217.710 ;
        RECT 33.245 217.060 33.505 217.450 ;
        RECT 33.675 217.230 33.955 217.710 ;
        RECT 31.765 216.470 32.115 217.040 ;
        RECT 32.350 216.890 34.000 217.060 ;
        RECT 32.285 216.550 33.425 216.720 ;
        RECT 32.285 216.300 32.455 216.550 ;
        RECT 33.595 216.380 34.000 216.890 ;
        RECT 34.185 216.960 35.395 217.710 ;
        RECT 34.185 216.420 34.705 216.960 ;
        RECT 35.625 216.890 35.835 217.710 ;
        RECT 36.005 216.910 36.335 217.540 ;
        RECT 31.425 216.130 32.455 216.300 ;
        RECT 33.245 216.210 34.000 216.380 ;
        RECT 34.875 216.250 35.395 216.790 ;
        RECT 36.005 216.310 36.255 216.910 ;
        RECT 36.505 216.890 36.735 217.710 ;
        RECT 36.945 217.210 37.245 217.540 ;
        RECT 37.415 217.230 37.690 217.710 ;
        RECT 36.425 216.470 36.755 216.720 ;
        RECT 31.425 215.330 31.735 216.130 ;
        RECT 33.245 215.960 33.505 216.210 ;
        RECT 31.905 215.160 32.215 215.960 ;
        RECT 32.385 215.790 33.505 215.960 ;
        RECT 32.385 215.330 32.645 215.790 ;
        RECT 32.815 215.160 33.070 215.620 ;
        RECT 33.245 215.330 33.505 215.790 ;
        RECT 33.675 215.160 33.960 216.030 ;
        RECT 34.185 215.160 35.395 216.250 ;
        RECT 35.625 215.160 35.835 216.300 ;
        RECT 36.005 215.330 36.335 216.310 ;
        RECT 36.945 216.300 37.115 217.210 ;
        RECT 37.870 217.060 38.165 217.450 ;
        RECT 38.335 217.230 38.590 217.710 ;
        RECT 38.765 217.060 39.025 217.450 ;
        RECT 39.195 217.230 39.475 217.710 ;
        RECT 37.285 216.470 37.635 217.040 ;
        RECT 37.870 216.890 39.520 217.060 ;
        RECT 39.705 216.985 39.995 217.710 ;
        RECT 37.805 216.550 38.945 216.720 ;
        RECT 37.805 216.300 37.975 216.550 ;
        RECT 39.115 216.380 39.520 216.890 ;
        RECT 36.505 215.160 36.735 216.300 ;
        RECT 36.945 216.130 37.975 216.300 ;
        RECT 38.765 216.210 39.520 216.380 ;
        RECT 40.170 216.970 40.425 217.540 ;
        RECT 40.595 217.310 40.925 217.710 ;
        RECT 41.350 217.175 41.880 217.540 ;
        RECT 41.350 217.140 41.525 217.175 ;
        RECT 40.595 216.970 41.525 217.140 ;
        RECT 36.945 215.330 37.255 216.130 ;
        RECT 38.765 215.960 39.025 216.210 ;
        RECT 37.425 215.160 37.735 215.960 ;
        RECT 37.905 215.790 39.025 215.960 ;
        RECT 37.905 215.330 38.165 215.790 ;
        RECT 38.335 215.160 38.590 215.620 ;
        RECT 38.765 215.330 39.025 215.790 ;
        RECT 39.195 215.160 39.480 216.030 ;
        RECT 39.705 215.160 39.995 216.325 ;
        RECT 40.170 216.300 40.340 216.970 ;
        RECT 40.595 216.800 40.765 216.970 ;
        RECT 40.510 216.470 40.765 216.800 ;
        RECT 40.990 216.470 41.185 216.800 ;
        RECT 40.170 215.330 40.505 216.300 ;
        RECT 40.675 215.160 40.845 216.300 ;
        RECT 41.015 215.500 41.185 216.470 ;
        RECT 41.355 215.840 41.525 216.970 ;
        RECT 41.695 216.180 41.865 216.980 ;
        RECT 42.070 216.690 42.345 217.540 ;
        RECT 42.065 216.520 42.345 216.690 ;
        RECT 42.070 216.380 42.345 216.520 ;
        RECT 42.515 216.180 42.705 217.540 ;
        RECT 42.885 217.175 43.395 217.710 ;
        RECT 43.615 216.900 43.860 217.505 ;
        RECT 44.310 216.970 44.565 217.540 ;
        RECT 44.735 217.310 45.065 217.710 ;
        RECT 45.490 217.175 46.020 217.540 ;
        RECT 45.490 217.140 45.665 217.175 ;
        RECT 44.735 216.970 45.665 217.140 ;
        RECT 46.210 217.030 46.485 217.540 ;
        RECT 42.905 216.730 44.135 216.900 ;
        RECT 41.695 216.010 42.705 216.180 ;
        RECT 42.875 216.165 43.625 216.355 ;
        RECT 41.355 215.670 42.480 215.840 ;
        RECT 42.875 215.500 43.045 216.165 ;
        RECT 43.795 215.920 44.135 216.730 ;
        RECT 41.015 215.330 43.045 215.500 ;
        RECT 43.215 215.160 43.385 215.920 ;
        RECT 43.620 215.510 44.135 215.920 ;
        RECT 44.310 216.300 44.480 216.970 ;
        RECT 44.735 216.800 44.905 216.970 ;
        RECT 44.650 216.470 44.905 216.800 ;
        RECT 45.130 216.470 45.325 216.800 ;
        RECT 44.310 215.330 44.645 216.300 ;
        RECT 44.815 215.160 44.985 216.300 ;
        RECT 45.155 215.500 45.325 216.470 ;
        RECT 45.495 215.840 45.665 216.970 ;
        RECT 45.835 216.180 46.005 216.980 ;
        RECT 46.205 216.860 46.485 217.030 ;
        RECT 46.210 216.380 46.485 216.860 ;
        RECT 46.655 216.180 46.845 217.540 ;
        RECT 47.025 217.175 47.535 217.710 ;
        RECT 47.755 216.900 48.000 217.505 ;
        RECT 47.045 216.730 48.275 216.900 ;
        RECT 48.505 216.890 48.715 217.710 ;
        RECT 48.885 216.910 49.215 217.540 ;
        RECT 45.835 216.010 46.845 216.180 ;
        RECT 47.015 216.165 47.765 216.355 ;
        RECT 45.495 215.670 46.620 215.840 ;
        RECT 47.015 215.500 47.185 216.165 ;
        RECT 47.935 215.920 48.275 216.730 ;
        RECT 48.885 216.310 49.135 216.910 ;
        RECT 49.385 216.890 49.615 217.710 ;
        RECT 49.825 217.210 50.125 217.540 ;
        RECT 50.295 217.230 50.570 217.710 ;
        RECT 49.305 216.470 49.635 216.720 ;
        RECT 45.155 215.330 47.185 215.500 ;
        RECT 47.355 215.160 47.525 215.920 ;
        RECT 47.760 215.510 48.275 215.920 ;
        RECT 48.505 215.160 48.715 216.300 ;
        RECT 48.885 215.330 49.215 216.310 ;
        RECT 49.825 216.300 49.995 217.210 ;
        RECT 50.750 217.060 51.045 217.450 ;
        RECT 51.215 217.230 51.470 217.710 ;
        RECT 51.645 217.060 51.905 217.450 ;
        RECT 52.075 217.230 52.355 217.710 ;
        RECT 50.165 216.470 50.515 217.040 ;
        RECT 50.750 216.890 52.400 217.060 ;
        RECT 52.585 216.985 52.875 217.710 ;
        RECT 50.685 216.550 51.825 216.720 ;
        RECT 50.685 216.300 50.855 216.550 ;
        RECT 51.995 216.380 52.400 216.890 ;
        RECT 49.385 215.160 49.615 216.300 ;
        RECT 49.825 216.130 50.855 216.300 ;
        RECT 51.645 216.210 52.400 216.380 ;
        RECT 53.050 216.970 53.305 217.540 ;
        RECT 53.475 217.310 53.805 217.710 ;
        RECT 54.230 217.175 54.760 217.540 ;
        RECT 54.230 217.140 54.405 217.175 ;
        RECT 53.475 216.970 54.405 217.140 ;
        RECT 49.825 215.330 50.135 216.130 ;
        RECT 51.645 215.960 51.905 216.210 ;
        RECT 50.305 215.160 50.615 215.960 ;
        RECT 50.785 215.790 51.905 215.960 ;
        RECT 50.785 215.330 51.045 215.790 ;
        RECT 51.215 215.160 51.470 215.620 ;
        RECT 51.645 215.330 51.905 215.790 ;
        RECT 52.075 215.160 52.360 216.030 ;
        RECT 52.585 215.160 52.875 216.325 ;
        RECT 53.050 216.300 53.220 216.970 ;
        RECT 53.475 216.800 53.645 216.970 ;
        RECT 53.390 216.470 53.645 216.800 ;
        RECT 53.870 216.470 54.065 216.800 ;
        RECT 53.050 215.330 53.385 216.300 ;
        RECT 53.555 215.160 53.725 216.300 ;
        RECT 53.895 215.500 54.065 216.470 ;
        RECT 54.235 215.840 54.405 216.970 ;
        RECT 54.575 216.180 54.745 216.980 ;
        RECT 54.950 216.690 55.225 217.540 ;
        RECT 54.945 216.520 55.225 216.690 ;
        RECT 54.950 216.380 55.225 216.520 ;
        RECT 55.395 216.180 55.585 217.540 ;
        RECT 55.765 217.175 56.275 217.710 ;
        RECT 56.495 216.900 56.740 217.505 ;
        RECT 57.185 216.960 58.395 217.710 ;
        RECT 58.625 217.230 58.905 217.710 ;
        RECT 59.075 217.060 59.335 217.450 ;
        RECT 59.510 217.230 59.765 217.710 ;
        RECT 59.935 217.060 60.230 217.450 ;
        RECT 60.410 217.230 60.685 217.710 ;
        RECT 60.855 217.210 61.155 217.540 ;
        RECT 55.785 216.730 57.015 216.900 ;
        RECT 54.575 216.010 55.585 216.180 ;
        RECT 55.755 216.165 56.505 216.355 ;
        RECT 54.235 215.670 55.360 215.840 ;
        RECT 55.755 215.500 55.925 216.165 ;
        RECT 56.675 215.920 57.015 216.730 ;
        RECT 57.185 216.420 57.705 216.960 ;
        RECT 58.580 216.890 60.230 217.060 ;
        RECT 57.875 216.250 58.395 216.790 ;
        RECT 53.895 215.330 55.925 215.500 ;
        RECT 56.095 215.160 56.265 215.920 ;
        RECT 56.500 215.510 57.015 215.920 ;
        RECT 57.185 215.160 58.395 216.250 ;
        RECT 58.580 216.380 58.985 216.890 ;
        RECT 59.155 216.550 60.295 216.720 ;
        RECT 58.580 216.210 59.335 216.380 ;
        RECT 58.620 215.160 58.905 216.030 ;
        RECT 59.075 215.960 59.335 216.210 ;
        RECT 60.125 216.300 60.295 216.550 ;
        RECT 60.465 216.470 60.815 217.040 ;
        RECT 60.985 216.300 61.155 217.210 ;
        RECT 62.305 216.890 62.515 217.710 ;
        RECT 62.685 216.910 63.015 217.540 ;
        RECT 62.685 216.310 62.935 216.910 ;
        RECT 63.185 216.890 63.415 217.710 ;
        RECT 63.665 216.890 63.895 217.710 ;
        RECT 64.065 216.910 64.395 217.540 ;
        RECT 63.105 216.470 63.435 216.720 ;
        RECT 63.645 216.470 63.975 216.720 ;
        RECT 64.145 216.310 64.395 216.910 ;
        RECT 64.565 216.890 64.775 217.710 ;
        RECT 65.465 216.985 65.755 217.710 ;
        RECT 65.925 217.210 66.225 217.540 ;
        RECT 66.395 217.230 66.670 217.710 ;
        RECT 60.125 216.130 61.155 216.300 ;
        RECT 59.075 215.790 60.195 215.960 ;
        RECT 59.075 215.330 59.335 215.790 ;
        RECT 59.510 215.160 59.765 215.620 ;
        RECT 59.935 215.330 60.195 215.790 ;
        RECT 60.365 215.160 60.675 215.960 ;
        RECT 60.845 215.330 61.155 216.130 ;
        RECT 62.305 215.160 62.515 216.300 ;
        RECT 62.685 215.330 63.015 216.310 ;
        RECT 63.185 215.160 63.415 216.300 ;
        RECT 63.665 215.160 63.895 216.300 ;
        RECT 64.065 215.330 64.395 216.310 ;
        RECT 64.565 215.160 64.775 216.300 ;
        RECT 65.465 215.160 65.755 216.325 ;
        RECT 65.925 216.300 66.095 217.210 ;
        RECT 66.850 217.060 67.145 217.450 ;
        RECT 67.315 217.230 67.570 217.710 ;
        RECT 67.745 217.060 68.005 217.450 ;
        RECT 68.175 217.230 68.455 217.710 ;
        RECT 69.345 217.080 69.675 217.440 ;
        RECT 70.295 217.250 70.545 217.710 ;
        RECT 70.715 217.250 71.275 217.540 ;
        RECT 66.265 216.470 66.615 217.040 ;
        RECT 66.850 216.890 68.500 217.060 ;
        RECT 69.345 216.890 70.735 217.080 ;
        RECT 66.785 216.550 67.925 216.720 ;
        RECT 66.785 216.300 66.955 216.550 ;
        RECT 68.095 216.380 68.500 216.890 ;
        RECT 70.565 216.800 70.735 216.890 ;
        RECT 65.925 216.130 66.955 216.300 ;
        RECT 67.745 216.210 68.500 216.380 ;
        RECT 69.160 216.470 69.835 216.720 ;
        RECT 70.055 216.470 70.395 216.720 ;
        RECT 70.565 216.470 70.855 216.800 ;
        RECT 65.925 215.330 66.235 216.130 ;
        RECT 67.745 215.960 68.005 216.210 ;
        RECT 69.160 216.110 69.425 216.470 ;
        RECT 70.565 216.220 70.735 216.470 ;
        RECT 69.795 216.050 70.735 216.220 ;
        RECT 66.405 215.160 66.715 215.960 ;
        RECT 66.885 215.790 68.005 215.960 ;
        RECT 66.885 215.330 67.145 215.790 ;
        RECT 67.315 215.160 67.570 215.620 ;
        RECT 67.745 215.330 68.005 215.790 ;
        RECT 68.175 215.160 68.460 216.030 ;
        RECT 69.345 215.160 69.625 215.830 ;
        RECT 69.795 215.500 70.095 216.050 ;
        RECT 71.025 215.880 71.275 217.250 ;
        RECT 71.445 216.940 74.955 217.710 ;
        RECT 75.125 217.210 75.425 217.540 ;
        RECT 75.595 217.230 75.870 217.710 ;
        RECT 71.445 216.420 73.095 216.940 ;
        RECT 73.265 216.250 74.955 216.770 ;
        RECT 70.295 215.160 70.625 215.880 ;
        RECT 70.815 215.330 71.275 215.880 ;
        RECT 71.445 215.160 74.955 216.250 ;
        RECT 75.125 216.300 75.295 217.210 ;
        RECT 76.050 217.060 76.345 217.450 ;
        RECT 76.515 217.230 76.770 217.710 ;
        RECT 76.945 217.060 77.205 217.450 ;
        RECT 77.375 217.230 77.655 217.710 ;
        RECT 75.465 216.470 75.815 217.040 ;
        RECT 76.050 216.890 77.700 217.060 ;
        RECT 78.345 216.985 78.635 217.710 ;
        RECT 78.805 217.250 79.365 217.540 ;
        RECT 79.535 217.250 79.785 217.710 ;
        RECT 75.985 216.550 77.125 216.720 ;
        RECT 75.985 216.300 76.155 216.550 ;
        RECT 77.295 216.380 77.700 216.890 ;
        RECT 75.125 216.130 76.155 216.300 ;
        RECT 76.945 216.210 77.700 216.380 ;
        RECT 75.125 215.330 75.435 216.130 ;
        RECT 76.945 215.960 77.205 216.210 ;
        RECT 75.605 215.160 75.915 215.960 ;
        RECT 76.085 215.790 77.205 215.960 ;
        RECT 76.085 215.330 76.345 215.790 ;
        RECT 76.515 215.160 76.770 215.620 ;
        RECT 76.945 215.330 77.205 215.790 ;
        RECT 77.375 215.160 77.660 216.030 ;
        RECT 78.345 215.160 78.635 216.325 ;
        RECT 78.805 215.880 79.055 217.250 ;
        RECT 80.405 217.080 80.735 217.440 ;
        RECT 79.345 216.890 80.735 217.080 ;
        RECT 81.105 216.940 84.615 217.710 ;
        RECT 84.985 217.080 85.315 217.440 ;
        RECT 85.935 217.250 86.185 217.710 ;
        RECT 86.355 217.250 86.915 217.540 ;
        RECT 79.345 216.800 79.515 216.890 ;
        RECT 79.225 216.470 79.515 216.800 ;
        RECT 79.685 216.470 80.025 216.720 ;
        RECT 80.245 216.470 80.920 216.720 ;
        RECT 79.345 216.220 79.515 216.470 ;
        RECT 79.345 216.050 80.285 216.220 ;
        RECT 80.655 216.110 80.920 216.470 ;
        RECT 81.105 216.420 82.755 216.940 ;
        RECT 84.985 216.890 86.375 217.080 ;
        RECT 86.205 216.800 86.375 216.890 ;
        RECT 82.925 216.250 84.615 216.770 ;
        RECT 78.805 215.330 79.265 215.880 ;
        RECT 79.455 215.160 79.785 215.880 ;
        RECT 79.985 215.500 80.285 216.050 ;
        RECT 80.455 215.160 80.735 215.830 ;
        RECT 81.105 215.160 84.615 216.250 ;
        RECT 84.800 216.470 85.475 216.720 ;
        RECT 85.695 216.470 86.035 216.720 ;
        RECT 86.205 216.470 86.495 216.800 ;
        RECT 84.800 216.110 85.065 216.470 ;
        RECT 86.205 216.220 86.375 216.470 ;
        RECT 85.435 216.050 86.375 216.220 ;
        RECT 84.985 215.160 85.265 215.830 ;
        RECT 85.435 215.500 85.735 216.050 ;
        RECT 86.665 215.880 86.915 217.250 ;
        RECT 85.935 215.160 86.265 215.880 ;
        RECT 86.455 215.330 86.915 215.880 ;
        RECT 87.085 217.210 87.385 217.540 ;
        RECT 87.555 217.230 87.830 217.710 ;
        RECT 87.085 216.300 87.255 217.210 ;
        RECT 88.010 217.060 88.305 217.450 ;
        RECT 88.475 217.230 88.730 217.710 ;
        RECT 88.905 217.060 89.165 217.450 ;
        RECT 89.335 217.230 89.615 217.710 ;
        RECT 87.425 216.470 87.775 217.040 ;
        RECT 88.010 216.890 89.660 217.060 ;
        RECT 87.945 216.550 89.085 216.720 ;
        RECT 87.945 216.300 88.115 216.550 ;
        RECT 89.255 216.380 89.660 216.890 ;
        RECT 89.845 216.960 91.055 217.710 ;
        RECT 91.225 216.985 91.515 217.710 ;
        RECT 89.845 216.420 90.365 216.960 ;
        RECT 91.685 216.940 94.275 217.710 ;
        RECT 87.085 216.130 88.115 216.300 ;
        RECT 88.905 216.210 89.660 216.380 ;
        RECT 90.535 216.250 91.055 216.790 ;
        RECT 91.685 216.420 92.895 216.940 ;
        RECT 94.965 216.890 95.175 217.710 ;
        RECT 95.345 216.910 95.675 217.540 ;
        RECT 87.085 215.330 87.395 216.130 ;
        RECT 88.905 215.960 89.165 216.210 ;
        RECT 87.565 215.160 87.875 215.960 ;
        RECT 88.045 215.790 89.165 215.960 ;
        RECT 88.045 215.330 88.305 215.790 ;
        RECT 88.475 215.160 88.730 215.620 ;
        RECT 88.905 215.330 89.165 215.790 ;
        RECT 89.335 215.160 89.620 216.030 ;
        RECT 89.845 215.160 91.055 216.250 ;
        RECT 91.225 215.160 91.515 216.325 ;
        RECT 93.065 216.250 94.275 216.770 ;
        RECT 95.345 216.310 95.595 216.910 ;
        RECT 95.845 216.890 96.075 217.710 ;
        RECT 96.285 216.970 96.545 217.710 ;
        RECT 96.795 216.890 96.985 217.360 ;
        RECT 97.235 217.210 97.485 217.710 ;
        RECT 97.815 217.140 97.985 217.490 ;
        RECT 98.185 217.310 98.515 217.710 ;
        RECT 98.685 217.140 98.855 217.490 ;
        RECT 99.075 217.310 99.455 217.710 ;
        RECT 96.815 216.800 96.985 216.890 ;
        RECT 97.655 216.970 99.465 217.140 ;
        RECT 95.765 216.470 96.095 216.720 ;
        RECT 91.685 215.160 94.275 216.250 ;
        RECT 94.965 215.160 95.175 216.300 ;
        RECT 95.345 215.330 95.675 216.310 ;
        RECT 95.845 215.160 96.075 216.300 ;
        RECT 96.305 215.840 96.645 216.800 ;
        RECT 96.815 216.470 97.415 216.800 ;
        RECT 96.815 215.730 96.985 216.470 ;
        RECT 97.655 216.220 97.825 216.970 ;
        RECT 96.285 215.160 96.565 215.660 ;
        RECT 96.795 215.340 96.985 215.730 ;
        RECT 97.235 216.050 97.825 216.220 ;
        RECT 97.995 216.175 98.165 216.800 ;
        RECT 98.395 216.345 98.725 216.800 ;
        RECT 97.235 215.345 97.565 216.050 ;
        RECT 97.995 215.420 98.355 216.175 ;
        RECT 98.535 216.010 98.725 216.345 ;
        RECT 98.955 216.350 99.125 216.800 ;
        RECT 99.295 216.720 99.465 216.970 ;
        RECT 99.635 217.070 99.885 217.540 ;
        RECT 100.055 217.240 100.225 217.710 ;
        RECT 100.395 217.070 100.725 217.540 ;
        RECT 100.895 217.240 101.065 217.710 ;
        RECT 101.435 217.160 101.605 217.540 ;
        RECT 101.785 217.330 102.115 217.710 ;
        RECT 99.635 216.890 101.165 217.070 ;
        RECT 101.435 216.990 102.100 217.160 ;
        RECT 102.295 217.035 102.555 217.540 ;
        RECT 99.295 216.550 100.755 216.720 ;
        RECT 98.955 216.180 99.390 216.350 ;
        RECT 100.925 216.340 101.165 216.890 ;
        RECT 101.365 216.440 101.705 216.810 ;
        RECT 101.930 216.735 102.100 216.990 ;
        RECT 99.595 216.170 101.165 216.340 ;
        RECT 101.930 216.405 102.205 216.735 ;
        RECT 101.930 216.260 102.100 216.405 ;
        RECT 98.535 215.420 98.835 216.010 ;
        RECT 99.120 215.160 99.370 216.000 ;
        RECT 99.595 215.330 99.845 216.170 ;
        RECT 100.015 215.160 100.265 216.000 ;
        RECT 100.435 215.330 100.685 216.170 ;
        RECT 101.425 216.090 102.100 216.260 ;
        RECT 102.375 216.235 102.555 217.035 ;
        RECT 102.725 216.960 103.935 217.710 ;
        RECT 104.105 216.985 104.395 217.710 ;
        RECT 104.655 217.160 104.825 217.540 ;
        RECT 105.040 217.330 105.370 217.710 ;
        RECT 104.655 216.990 105.370 217.160 ;
        RECT 102.725 216.420 103.245 216.960 ;
        RECT 103.415 216.250 103.935 216.790 ;
        RECT 104.565 216.440 104.920 216.810 ;
        RECT 105.200 216.800 105.370 216.990 ;
        RECT 105.540 216.965 105.795 217.540 ;
        RECT 105.200 216.470 105.455 216.800 ;
        RECT 100.855 215.160 101.105 216.000 ;
        RECT 101.425 215.330 101.605 216.090 ;
        RECT 101.785 215.160 102.115 215.920 ;
        RECT 102.285 215.330 102.555 216.235 ;
        RECT 102.725 215.160 103.935 216.250 ;
        RECT 104.105 215.160 104.395 216.325 ;
        RECT 105.200 216.260 105.370 216.470 ;
        RECT 104.655 216.090 105.370 216.260 ;
        RECT 105.625 216.235 105.795 216.965 ;
        RECT 105.970 216.870 106.230 217.710 ;
        RECT 107.330 217.160 107.585 217.450 ;
        RECT 107.755 217.330 108.085 217.710 ;
        RECT 107.330 216.990 108.080 217.160 ;
        RECT 104.655 215.330 104.825 216.090 ;
        RECT 105.040 215.160 105.370 215.920 ;
        RECT 105.540 215.330 105.795 216.235 ;
        RECT 105.970 215.160 106.230 216.310 ;
        RECT 107.330 216.170 107.680 216.820 ;
        RECT 107.850 216.000 108.080 216.990 ;
        RECT 107.330 215.830 108.080 216.000 ;
        RECT 107.330 215.330 107.585 215.830 ;
        RECT 107.755 215.160 108.085 215.660 ;
        RECT 108.255 215.330 108.425 217.450 ;
        RECT 108.785 217.350 109.115 217.710 ;
        RECT 109.285 217.320 109.780 217.490 ;
        RECT 109.985 217.320 110.840 217.490 ;
        RECT 108.655 216.130 109.115 217.180 ;
        RECT 108.595 215.345 108.920 216.130 ;
        RECT 109.285 215.960 109.455 217.320 ;
        RECT 109.625 216.410 109.975 217.030 ;
        RECT 110.145 216.810 110.500 217.030 ;
        RECT 110.145 216.220 110.315 216.810 ;
        RECT 110.670 216.610 110.840 217.320 ;
        RECT 111.715 217.250 112.045 217.710 ;
        RECT 112.255 217.350 112.605 217.520 ;
        RECT 111.045 216.780 111.835 217.030 ;
        RECT 112.255 216.960 112.515 217.350 ;
        RECT 112.825 217.260 113.775 217.540 ;
        RECT 113.945 217.270 114.135 217.710 ;
        RECT 114.305 217.330 115.375 217.500 ;
        RECT 112.005 216.610 112.175 216.790 ;
        RECT 109.285 215.790 109.680 215.960 ;
        RECT 109.850 215.830 110.315 216.220 ;
        RECT 110.485 216.440 112.175 216.610 ;
        RECT 109.510 215.660 109.680 215.790 ;
        RECT 110.485 215.660 110.655 216.440 ;
        RECT 112.345 216.270 112.515 216.960 ;
        RECT 111.015 216.100 112.515 216.270 ;
        RECT 112.705 216.300 112.915 217.090 ;
        RECT 113.085 216.470 113.435 217.090 ;
        RECT 113.605 216.480 113.775 217.260 ;
        RECT 114.305 217.100 114.475 217.330 ;
        RECT 113.945 216.930 114.475 217.100 ;
        RECT 113.945 216.650 114.165 216.930 ;
        RECT 114.645 216.760 114.885 217.160 ;
        RECT 113.605 216.310 114.010 216.480 ;
        RECT 114.345 216.390 114.885 216.760 ;
        RECT 115.055 216.975 115.375 217.330 ;
        RECT 115.620 217.250 115.925 217.710 ;
        RECT 116.095 217.000 116.345 217.530 ;
        RECT 115.055 216.800 115.380 216.975 ;
        RECT 115.055 216.500 115.970 216.800 ;
        RECT 115.230 216.470 115.970 216.500 ;
        RECT 112.705 216.140 113.380 216.300 ;
        RECT 113.840 216.220 114.010 216.310 ;
        RECT 112.705 216.130 113.670 216.140 ;
        RECT 112.345 215.960 112.515 216.100 ;
        RECT 109.090 215.160 109.340 215.620 ;
        RECT 109.510 215.330 109.760 215.660 ;
        RECT 109.975 215.330 110.655 215.660 ;
        RECT 110.825 215.760 111.900 215.930 ;
        RECT 112.345 215.790 112.905 215.960 ;
        RECT 113.210 215.840 113.670 216.130 ;
        RECT 113.840 216.050 115.060 216.220 ;
        RECT 110.825 215.420 110.995 215.760 ;
        RECT 111.230 215.160 111.560 215.590 ;
        RECT 111.730 215.420 111.900 215.760 ;
        RECT 112.195 215.160 112.565 215.620 ;
        RECT 112.735 215.330 112.905 215.790 ;
        RECT 113.840 215.670 114.010 216.050 ;
        RECT 115.230 215.880 115.400 216.470 ;
        RECT 116.140 216.350 116.345 217.000 ;
        RECT 116.515 216.955 116.765 217.710 ;
        RECT 116.985 216.985 117.275 217.710 ;
        RECT 117.505 217.230 117.785 217.710 ;
        RECT 117.955 217.060 118.215 217.450 ;
        RECT 118.390 217.230 118.645 217.710 ;
        RECT 118.815 217.060 119.110 217.450 ;
        RECT 119.290 217.230 119.565 217.710 ;
        RECT 119.735 217.210 120.035 217.540 ;
        RECT 120.265 217.230 120.545 217.710 ;
        RECT 113.140 215.330 114.010 215.670 ;
        RECT 114.600 215.710 115.400 215.880 ;
        RECT 114.180 215.160 114.430 215.620 ;
        RECT 114.600 215.420 114.770 215.710 ;
        RECT 114.950 215.160 115.280 215.540 ;
        RECT 115.620 215.160 115.925 216.300 ;
        RECT 116.095 215.470 116.345 216.350 ;
        RECT 117.460 216.890 119.110 217.060 ;
        RECT 117.460 216.380 117.865 216.890 ;
        RECT 118.035 216.550 119.175 216.720 ;
        RECT 116.515 215.160 116.765 216.300 ;
        RECT 116.985 215.160 117.275 216.325 ;
        RECT 117.460 216.210 118.215 216.380 ;
        RECT 117.500 215.160 117.785 216.030 ;
        RECT 117.955 215.960 118.215 216.210 ;
        RECT 119.005 216.300 119.175 216.550 ;
        RECT 119.345 216.470 119.695 217.040 ;
        RECT 119.865 216.300 120.035 217.210 ;
        RECT 120.715 217.060 120.975 217.450 ;
        RECT 121.150 217.230 121.405 217.710 ;
        RECT 121.575 217.060 121.870 217.450 ;
        RECT 122.050 217.230 122.325 217.710 ;
        RECT 122.495 217.210 122.795 217.540 ;
        RECT 119.005 216.130 120.035 216.300 ;
        RECT 120.220 216.890 121.870 217.060 ;
        RECT 120.220 216.380 120.625 216.890 ;
        RECT 120.795 216.550 121.935 216.720 ;
        RECT 120.220 216.210 120.975 216.380 ;
        RECT 117.955 215.790 119.075 215.960 ;
        RECT 117.955 215.330 118.215 215.790 ;
        RECT 118.390 215.160 118.645 215.620 ;
        RECT 118.815 215.330 119.075 215.790 ;
        RECT 119.245 215.160 119.555 215.960 ;
        RECT 119.725 215.330 120.035 216.130 ;
        RECT 120.260 215.160 120.545 216.030 ;
        RECT 120.715 215.960 120.975 216.210 ;
        RECT 121.765 216.300 121.935 216.550 ;
        RECT 122.105 216.470 122.455 217.040 ;
        RECT 122.625 216.300 122.795 217.210 ;
        RECT 123.430 216.870 123.690 217.710 ;
        RECT 123.865 216.965 124.120 217.540 ;
        RECT 124.290 217.330 124.620 217.710 ;
        RECT 124.835 217.160 125.005 217.540 ;
        RECT 124.290 216.990 125.005 217.160 ;
        RECT 126.230 217.250 126.980 217.540 ;
        RECT 127.490 217.250 127.820 217.710 ;
        RECT 121.765 216.130 122.795 216.300 ;
        RECT 120.715 215.790 121.835 215.960 ;
        RECT 120.715 215.330 120.975 215.790 ;
        RECT 121.150 215.160 121.405 215.620 ;
        RECT 121.575 215.330 121.835 215.790 ;
        RECT 122.005 215.160 122.315 215.960 ;
        RECT 122.485 215.330 122.795 216.130 ;
        RECT 123.430 215.160 123.690 216.310 ;
        RECT 123.865 216.235 124.035 216.965 ;
        RECT 124.290 216.800 124.460 216.990 ;
        RECT 124.205 216.470 124.460 216.800 ;
        RECT 124.290 216.260 124.460 216.470 ;
        RECT 124.740 216.440 125.095 216.810 ;
        RECT 123.865 215.330 124.120 216.235 ;
        RECT 124.290 216.090 125.005 216.260 ;
        RECT 124.290 215.160 124.620 215.920 ;
        RECT 124.835 215.330 125.005 216.090 ;
        RECT 126.230 215.960 126.600 217.250 ;
        RECT 128.040 217.060 128.310 217.270 ;
        RECT 126.975 216.890 128.310 217.060 ;
        RECT 128.485 217.035 128.745 217.540 ;
        RECT 128.925 217.330 129.255 217.710 ;
        RECT 129.435 217.160 129.605 217.540 ;
        RECT 126.975 216.720 127.145 216.890 ;
        RECT 126.770 216.470 127.145 216.720 ;
        RECT 127.315 216.480 127.790 216.720 ;
        RECT 127.960 216.480 128.310 216.720 ;
        RECT 126.975 216.300 127.145 216.470 ;
        RECT 126.975 216.130 128.310 216.300 ;
        RECT 128.030 215.970 128.310 216.130 ;
        RECT 128.485 216.235 128.655 217.035 ;
        RECT 128.940 216.990 129.605 217.160 ;
        RECT 128.940 216.735 129.110 216.990 ;
        RECT 129.865 216.985 130.155 217.710 ;
        RECT 130.325 216.940 133.835 217.710 ;
        RECT 134.005 216.970 134.265 217.540 ;
        RECT 134.435 217.310 134.820 217.710 ;
        RECT 134.990 217.140 135.245 217.540 ;
        RECT 134.435 216.970 135.245 217.140 ;
        RECT 135.435 216.970 135.680 217.540 ;
        RECT 135.850 217.310 136.235 217.710 ;
        RECT 136.405 217.140 136.660 217.540 ;
        RECT 135.850 216.970 136.660 217.140 ;
        RECT 136.850 216.970 137.275 217.540 ;
        RECT 137.445 217.310 137.830 217.710 ;
        RECT 138.000 217.140 138.435 217.540 ;
        RECT 137.445 216.970 138.435 217.140 ;
        RECT 138.605 217.035 138.865 217.540 ;
        RECT 139.045 217.330 139.375 217.710 ;
        RECT 139.555 217.160 139.725 217.540 ;
        RECT 128.825 216.405 129.110 216.735 ;
        RECT 129.345 216.440 129.675 216.810 ;
        RECT 130.325 216.420 131.975 216.940 ;
        RECT 128.940 216.260 129.110 216.405 ;
        RECT 126.230 215.790 127.400 215.960 ;
        RECT 126.685 215.160 126.900 215.620 ;
        RECT 127.070 215.330 127.400 215.790 ;
        RECT 127.570 215.160 127.820 215.960 ;
        RECT 128.485 215.330 128.755 216.235 ;
        RECT 128.940 216.090 129.605 216.260 ;
        RECT 128.925 215.160 129.255 215.920 ;
        RECT 129.435 215.330 129.605 216.090 ;
        RECT 129.865 215.160 130.155 216.325 ;
        RECT 132.145 216.250 133.835 216.770 ;
        RECT 130.325 215.160 133.835 216.250 ;
        RECT 134.005 216.300 134.190 216.970 ;
        RECT 134.435 216.800 134.785 216.970 ;
        RECT 135.435 216.800 135.605 216.970 ;
        RECT 135.850 216.800 136.200 216.970 ;
        RECT 136.850 216.800 137.200 216.970 ;
        RECT 137.445 216.800 137.780 216.970 ;
        RECT 134.360 216.470 134.785 216.800 ;
        RECT 134.005 215.330 134.265 216.300 ;
        RECT 134.435 215.950 134.785 216.470 ;
        RECT 134.955 216.300 135.605 216.800 ;
        RECT 135.775 216.470 136.200 216.800 ;
        RECT 134.955 216.120 135.680 216.300 ;
        RECT 134.435 215.755 135.245 215.950 ;
        RECT 134.435 215.160 134.820 215.585 ;
        RECT 134.990 215.330 135.245 215.755 ;
        RECT 135.435 215.330 135.680 216.120 ;
        RECT 135.850 215.950 136.200 216.470 ;
        RECT 136.370 216.300 137.200 216.800 ;
        RECT 137.370 216.470 137.780 216.800 ;
        RECT 136.370 216.120 137.275 216.300 ;
        RECT 135.850 215.755 136.680 215.950 ;
        RECT 135.850 215.160 136.235 215.585 ;
        RECT 136.405 215.330 136.680 215.755 ;
        RECT 136.850 215.330 137.275 216.120 ;
        RECT 137.445 215.925 137.780 216.470 ;
        RECT 137.950 216.095 138.435 216.800 ;
        RECT 138.605 216.235 138.775 217.035 ;
        RECT 139.060 216.990 139.725 217.160 ;
        RECT 140.995 217.160 141.165 217.540 ;
        RECT 141.380 217.330 141.710 217.710 ;
        RECT 140.995 216.990 141.710 217.160 ;
        RECT 139.060 216.735 139.230 216.990 ;
        RECT 138.945 216.405 139.230 216.735 ;
        RECT 139.465 216.440 139.795 216.810 ;
        RECT 140.905 216.440 141.260 216.810 ;
        RECT 141.540 216.800 141.710 216.990 ;
        RECT 141.880 216.965 142.135 217.540 ;
        RECT 141.540 216.470 141.795 216.800 ;
        RECT 139.060 216.260 139.230 216.405 ;
        RECT 141.540 216.260 141.710 216.470 ;
        RECT 137.445 215.755 138.435 215.925 ;
        RECT 137.445 215.160 137.830 215.585 ;
        RECT 138.000 215.330 138.435 215.755 ;
        RECT 138.605 215.330 138.875 216.235 ;
        RECT 139.060 216.090 139.725 216.260 ;
        RECT 139.045 215.160 139.375 215.920 ;
        RECT 139.555 215.330 139.725 216.090 ;
        RECT 140.995 216.090 141.710 216.260 ;
        RECT 141.965 216.235 142.135 216.965 ;
        RECT 142.310 216.870 142.570 217.710 ;
        RECT 142.745 216.985 143.035 217.710 ;
        RECT 143.205 217.035 143.465 217.540 ;
        RECT 143.645 217.330 143.975 217.710 ;
        RECT 144.155 217.160 144.325 217.540 ;
        RECT 140.995 215.330 141.165 216.090 ;
        RECT 141.380 215.160 141.710 215.920 ;
        RECT 141.880 215.330 142.135 216.235 ;
        RECT 142.310 215.160 142.570 216.310 ;
        RECT 142.745 215.160 143.035 216.325 ;
        RECT 143.205 216.235 143.375 217.035 ;
        RECT 143.660 216.990 144.325 217.160 ;
        RECT 144.675 217.160 144.845 217.540 ;
        RECT 145.060 217.330 145.390 217.710 ;
        RECT 144.675 216.990 145.390 217.160 ;
        RECT 143.660 216.735 143.830 216.990 ;
        RECT 143.545 216.405 143.830 216.735 ;
        RECT 144.065 216.440 144.395 216.810 ;
        RECT 144.585 216.440 144.940 216.810 ;
        RECT 145.220 216.800 145.390 216.990 ;
        RECT 145.560 216.965 145.815 217.540 ;
        RECT 145.220 216.470 145.475 216.800 ;
        RECT 143.660 216.260 143.830 216.405 ;
        RECT 145.220 216.260 145.390 216.470 ;
        RECT 143.205 215.330 143.475 216.235 ;
        RECT 143.660 216.090 144.325 216.260 ;
        RECT 143.645 215.160 143.975 215.920 ;
        RECT 144.155 215.330 144.325 216.090 ;
        RECT 144.675 216.090 145.390 216.260 ;
        RECT 145.645 216.235 145.815 216.965 ;
        RECT 145.990 216.870 146.250 217.710 ;
        RECT 146.425 216.960 147.635 217.710 ;
        RECT 144.675 215.330 144.845 216.090 ;
        RECT 145.060 215.160 145.390 215.920 ;
        RECT 145.560 215.330 145.815 216.235 ;
        RECT 145.990 215.160 146.250 216.310 ;
        RECT 146.425 216.250 146.945 216.790 ;
        RECT 147.115 216.420 147.635 216.960 ;
        RECT 146.425 215.160 147.635 216.250 ;
        RECT 13.860 214.990 147.720 215.160 ;
        RECT 13.945 213.900 15.155 214.990 ;
        RECT 13.945 213.190 14.465 213.730 ;
        RECT 14.635 213.360 15.155 213.900 ;
        RECT 15.330 213.840 15.590 214.990 ;
        RECT 15.765 213.915 16.020 214.820 ;
        RECT 16.190 214.230 16.520 214.990 ;
        RECT 16.735 214.060 16.905 214.820 ;
        RECT 13.945 212.440 15.155 213.190 ;
        RECT 15.330 212.440 15.590 213.280 ;
        RECT 15.765 213.185 15.935 213.915 ;
        RECT 16.190 213.890 16.905 214.060 ;
        RECT 16.190 213.680 16.360 213.890 ;
        RECT 17.170 213.840 17.430 214.990 ;
        RECT 17.605 213.915 17.860 214.820 ;
        RECT 18.030 214.230 18.360 214.990 ;
        RECT 18.575 214.060 18.745 214.820 ;
        RECT 16.105 213.350 16.360 213.680 ;
        RECT 15.765 212.610 16.020 213.185 ;
        RECT 16.190 213.160 16.360 213.350 ;
        RECT 16.640 213.340 16.995 213.710 ;
        RECT 16.190 212.990 16.905 213.160 ;
        RECT 16.190 212.440 16.520 212.820 ;
        RECT 16.735 212.610 16.905 212.990 ;
        RECT 17.170 212.440 17.430 213.280 ;
        RECT 17.605 213.185 17.775 213.915 ;
        RECT 18.030 213.890 18.745 214.060 ;
        RECT 18.030 213.680 18.200 213.890 ;
        RECT 19.010 213.840 19.270 214.990 ;
        RECT 19.445 213.915 19.700 214.820 ;
        RECT 19.870 214.230 20.200 214.990 ;
        RECT 20.415 214.060 20.585 214.820 ;
        RECT 17.945 213.350 18.200 213.680 ;
        RECT 17.605 212.610 17.860 213.185 ;
        RECT 18.030 213.160 18.200 213.350 ;
        RECT 18.480 213.340 18.835 213.710 ;
        RECT 18.030 212.990 18.745 213.160 ;
        RECT 18.030 212.440 18.360 212.820 ;
        RECT 18.575 212.610 18.745 212.990 ;
        RECT 19.010 212.440 19.270 213.280 ;
        RECT 19.445 213.185 19.615 213.915 ;
        RECT 19.870 213.890 20.585 214.060 ;
        RECT 20.845 213.900 24.355 214.990 ;
        RECT 24.725 214.320 25.005 214.990 ;
        RECT 25.175 214.100 25.475 214.650 ;
        RECT 25.675 214.270 26.005 214.990 ;
        RECT 26.195 214.270 26.655 214.820 ;
        RECT 19.870 213.680 20.040 213.890 ;
        RECT 19.785 213.350 20.040 213.680 ;
        RECT 19.445 212.610 19.700 213.185 ;
        RECT 19.870 213.160 20.040 213.350 ;
        RECT 20.320 213.340 20.675 213.710 ;
        RECT 20.845 213.210 22.495 213.730 ;
        RECT 22.665 213.380 24.355 213.900 ;
        RECT 24.540 213.680 24.805 214.040 ;
        RECT 25.175 213.930 26.115 214.100 ;
        RECT 25.945 213.680 26.115 213.930 ;
        RECT 24.540 213.430 25.215 213.680 ;
        RECT 25.435 213.430 25.775 213.680 ;
        RECT 25.945 213.350 26.235 213.680 ;
        RECT 25.945 213.260 26.115 213.350 ;
        RECT 19.870 212.990 20.585 213.160 ;
        RECT 19.870 212.440 20.200 212.820 ;
        RECT 20.415 212.610 20.585 212.990 ;
        RECT 20.845 212.440 24.355 213.210 ;
        RECT 24.725 213.070 26.115 213.260 ;
        RECT 24.725 212.710 25.055 213.070 ;
        RECT 26.405 212.900 26.655 214.270 ;
        RECT 26.825 213.825 27.115 214.990 ;
        RECT 27.285 213.900 28.955 214.990 ;
        RECT 29.130 214.320 29.385 214.820 ;
        RECT 29.555 214.490 29.885 214.990 ;
        RECT 29.130 214.150 29.880 214.320 ;
        RECT 27.285 213.210 28.035 213.730 ;
        RECT 28.205 213.380 28.955 213.900 ;
        RECT 29.130 213.330 29.480 213.980 ;
        RECT 25.675 212.440 25.925 212.900 ;
        RECT 26.095 212.610 26.655 212.900 ;
        RECT 26.825 212.440 27.115 213.165 ;
        RECT 27.285 212.440 28.955 213.210 ;
        RECT 29.650 213.160 29.880 214.150 ;
        RECT 29.130 212.990 29.880 213.160 ;
        RECT 29.130 212.700 29.385 212.990 ;
        RECT 29.555 212.440 29.885 212.820 ;
        RECT 30.055 212.700 30.225 214.820 ;
        RECT 30.395 214.020 30.720 214.805 ;
        RECT 30.890 214.530 31.140 214.990 ;
        RECT 31.310 214.490 31.560 214.820 ;
        RECT 31.775 214.490 32.455 214.820 ;
        RECT 31.310 214.360 31.480 214.490 ;
        RECT 31.085 214.190 31.480 214.360 ;
        RECT 30.455 212.970 30.915 214.020 ;
        RECT 31.085 212.830 31.255 214.190 ;
        RECT 31.650 213.930 32.115 214.320 ;
        RECT 31.425 213.120 31.775 213.740 ;
        RECT 31.945 213.340 32.115 213.930 ;
        RECT 32.285 213.710 32.455 214.490 ;
        RECT 32.625 214.390 32.795 214.730 ;
        RECT 33.030 214.560 33.360 214.990 ;
        RECT 33.530 214.390 33.700 214.730 ;
        RECT 33.995 214.530 34.365 214.990 ;
        RECT 32.625 214.220 33.700 214.390 ;
        RECT 34.535 214.360 34.705 214.820 ;
        RECT 34.940 214.480 35.810 214.820 ;
        RECT 35.980 214.530 36.230 214.990 ;
        RECT 34.145 214.190 34.705 214.360 ;
        RECT 34.145 214.050 34.315 214.190 ;
        RECT 32.815 213.880 34.315 214.050 ;
        RECT 35.010 214.020 35.470 214.310 ;
        RECT 32.285 213.540 33.975 213.710 ;
        RECT 31.945 213.120 32.300 213.340 ;
        RECT 32.470 212.830 32.640 213.540 ;
        RECT 32.845 213.120 33.635 213.370 ;
        RECT 33.805 213.360 33.975 213.540 ;
        RECT 34.145 213.190 34.315 213.880 ;
        RECT 30.585 212.440 30.915 212.800 ;
        RECT 31.085 212.660 31.580 212.830 ;
        RECT 31.785 212.660 32.640 212.830 ;
        RECT 33.515 212.440 33.845 212.900 ;
        RECT 34.055 212.800 34.315 213.190 ;
        RECT 34.505 214.010 35.470 214.020 ;
        RECT 35.640 214.100 35.810 214.480 ;
        RECT 36.400 214.440 36.570 214.730 ;
        RECT 36.750 214.610 37.080 214.990 ;
        RECT 36.400 214.270 37.200 214.440 ;
        RECT 34.505 213.850 35.180 214.010 ;
        RECT 35.640 213.930 36.860 214.100 ;
        RECT 34.505 213.060 34.715 213.850 ;
        RECT 35.640 213.840 35.810 213.930 ;
        RECT 34.885 213.060 35.235 213.680 ;
        RECT 35.405 213.670 35.810 213.840 ;
        RECT 35.405 212.890 35.575 213.670 ;
        RECT 35.745 213.220 35.965 213.500 ;
        RECT 36.145 213.390 36.685 213.760 ;
        RECT 37.030 213.650 37.200 214.270 ;
        RECT 37.375 213.930 37.545 214.990 ;
        RECT 37.755 213.980 38.045 214.820 ;
        RECT 38.215 214.150 38.385 214.990 ;
        RECT 38.595 213.980 38.845 214.820 ;
        RECT 39.055 214.150 39.225 214.990 ;
        RECT 40.200 214.190 40.450 214.990 ;
        RECT 40.620 214.360 40.950 214.820 ;
        RECT 41.120 214.530 41.335 214.990 ;
        RECT 40.620 214.190 41.790 214.360 ;
        RECT 39.710 214.020 39.990 214.180 ;
        RECT 37.755 213.810 39.480 213.980 ;
        RECT 39.710 213.850 41.045 214.020 ;
        RECT 35.745 213.050 36.275 213.220 ;
        RECT 34.055 212.630 34.405 212.800 ;
        RECT 34.625 212.610 35.575 212.890 ;
        RECT 35.745 212.440 35.935 212.880 ;
        RECT 36.105 212.820 36.275 213.050 ;
        RECT 36.445 212.990 36.685 213.390 ;
        RECT 36.855 213.640 37.200 213.650 ;
        RECT 36.855 213.430 38.885 213.640 ;
        RECT 36.855 213.175 37.180 213.430 ;
        RECT 39.070 213.260 39.480 213.810 ;
        RECT 40.875 213.680 41.045 213.850 ;
        RECT 39.710 213.430 40.060 213.670 ;
        RECT 40.230 213.430 40.705 213.670 ;
        RECT 40.875 213.430 41.250 213.680 ;
        RECT 40.875 213.260 41.045 213.430 ;
        RECT 36.855 212.820 37.175 213.175 ;
        RECT 36.105 212.650 37.175 212.820 ;
        RECT 37.375 212.440 37.545 213.250 ;
        RECT 37.715 213.090 39.480 213.260 ;
        RECT 39.710 213.090 41.045 213.260 ;
        RECT 37.715 212.610 38.045 213.090 ;
        RECT 38.215 212.440 38.385 212.910 ;
        RECT 38.555 212.610 38.885 213.090 ;
        RECT 39.055 212.440 39.225 212.910 ;
        RECT 39.710 212.880 39.980 213.090 ;
        RECT 41.420 212.900 41.790 214.190 ;
        RECT 42.010 214.320 42.265 214.820 ;
        RECT 42.435 214.490 42.765 214.990 ;
        RECT 42.010 214.150 42.760 214.320 ;
        RECT 42.010 213.330 42.360 213.980 ;
        RECT 42.530 213.160 42.760 214.150 ;
        RECT 40.200 212.440 40.530 212.900 ;
        RECT 41.040 212.610 41.790 212.900 ;
        RECT 42.010 212.990 42.760 213.160 ;
        RECT 42.010 212.700 42.265 212.990 ;
        RECT 42.435 212.440 42.765 212.820 ;
        RECT 42.935 212.700 43.105 214.820 ;
        RECT 43.275 214.020 43.600 214.805 ;
        RECT 43.770 214.530 44.020 214.990 ;
        RECT 44.190 214.490 44.440 214.820 ;
        RECT 44.655 214.490 45.335 214.820 ;
        RECT 44.190 214.360 44.360 214.490 ;
        RECT 43.965 214.190 44.360 214.360 ;
        RECT 43.335 212.970 43.795 214.020 ;
        RECT 43.965 212.830 44.135 214.190 ;
        RECT 44.530 213.930 44.995 214.320 ;
        RECT 44.305 213.120 44.655 213.740 ;
        RECT 44.825 213.340 44.995 213.930 ;
        RECT 45.165 213.710 45.335 214.490 ;
        RECT 45.505 214.390 45.675 214.730 ;
        RECT 45.910 214.560 46.240 214.990 ;
        RECT 46.410 214.390 46.580 214.730 ;
        RECT 46.875 214.530 47.245 214.990 ;
        RECT 45.505 214.220 46.580 214.390 ;
        RECT 47.415 214.360 47.585 214.820 ;
        RECT 47.820 214.480 48.690 214.820 ;
        RECT 48.860 214.530 49.110 214.990 ;
        RECT 47.025 214.190 47.585 214.360 ;
        RECT 47.025 214.050 47.195 214.190 ;
        RECT 45.695 213.880 47.195 214.050 ;
        RECT 47.890 214.020 48.350 214.310 ;
        RECT 45.165 213.540 46.855 213.710 ;
        RECT 44.825 213.120 45.180 213.340 ;
        RECT 45.350 212.830 45.520 213.540 ;
        RECT 45.725 213.120 46.515 213.370 ;
        RECT 46.685 213.360 46.855 213.540 ;
        RECT 47.025 213.190 47.195 213.880 ;
        RECT 43.465 212.440 43.795 212.800 ;
        RECT 43.965 212.660 44.460 212.830 ;
        RECT 44.665 212.660 45.520 212.830 ;
        RECT 46.395 212.440 46.725 212.900 ;
        RECT 46.935 212.800 47.195 213.190 ;
        RECT 47.385 214.010 48.350 214.020 ;
        RECT 48.520 214.100 48.690 214.480 ;
        RECT 49.280 214.440 49.450 214.730 ;
        RECT 49.630 214.610 49.960 214.990 ;
        RECT 49.280 214.270 50.080 214.440 ;
        RECT 47.385 213.850 48.060 214.010 ;
        RECT 48.520 213.930 49.740 214.100 ;
        RECT 47.385 213.060 47.595 213.850 ;
        RECT 48.520 213.840 48.690 213.930 ;
        RECT 47.765 213.060 48.115 213.680 ;
        RECT 48.285 213.670 48.690 213.840 ;
        RECT 48.285 212.890 48.455 213.670 ;
        RECT 48.625 213.220 48.845 213.500 ;
        RECT 49.025 213.390 49.565 213.760 ;
        RECT 49.910 213.680 50.080 214.270 ;
        RECT 50.300 213.850 50.605 214.990 ;
        RECT 50.775 213.800 51.030 214.680 ;
        RECT 51.205 213.900 52.415 214.990 ;
        RECT 49.910 213.650 50.650 213.680 ;
        RECT 48.625 213.050 49.155 213.220 ;
        RECT 46.935 212.630 47.285 212.800 ;
        RECT 47.505 212.610 48.455 212.890 ;
        RECT 48.625 212.440 48.815 212.880 ;
        RECT 48.985 212.820 49.155 213.050 ;
        RECT 49.325 212.990 49.565 213.390 ;
        RECT 49.735 213.350 50.650 213.650 ;
        RECT 49.735 213.175 50.060 213.350 ;
        RECT 49.735 212.820 50.055 213.175 ;
        RECT 50.820 213.150 51.030 213.800 ;
        RECT 48.985 212.650 50.055 212.820 ;
        RECT 50.300 212.440 50.605 212.900 ;
        RECT 50.775 212.620 51.030 213.150 ;
        RECT 51.205 213.190 51.725 213.730 ;
        RECT 51.895 213.360 52.415 213.900 ;
        RECT 52.585 213.825 52.875 214.990 ;
        RECT 53.050 214.320 53.305 214.820 ;
        RECT 53.475 214.490 53.805 214.990 ;
        RECT 53.050 214.150 53.800 214.320 ;
        RECT 53.050 213.330 53.400 213.980 ;
        RECT 51.205 212.440 52.415 213.190 ;
        RECT 52.585 212.440 52.875 213.165 ;
        RECT 53.570 213.160 53.800 214.150 ;
        RECT 53.050 212.990 53.800 213.160 ;
        RECT 53.050 212.700 53.305 212.990 ;
        RECT 53.475 212.440 53.805 212.820 ;
        RECT 53.975 212.700 54.145 214.820 ;
        RECT 54.315 214.020 54.640 214.805 ;
        RECT 54.810 214.530 55.060 214.990 ;
        RECT 55.230 214.490 55.480 214.820 ;
        RECT 55.695 214.490 56.375 214.820 ;
        RECT 55.230 214.360 55.400 214.490 ;
        RECT 55.005 214.190 55.400 214.360 ;
        RECT 54.375 212.970 54.835 214.020 ;
        RECT 55.005 212.830 55.175 214.190 ;
        RECT 55.570 213.930 56.035 214.320 ;
        RECT 55.345 213.120 55.695 213.740 ;
        RECT 55.865 213.340 56.035 213.930 ;
        RECT 56.205 213.710 56.375 214.490 ;
        RECT 56.545 214.390 56.715 214.730 ;
        RECT 56.950 214.560 57.280 214.990 ;
        RECT 57.450 214.390 57.620 214.730 ;
        RECT 57.915 214.530 58.285 214.990 ;
        RECT 56.545 214.220 57.620 214.390 ;
        RECT 58.455 214.360 58.625 214.820 ;
        RECT 58.860 214.480 59.730 214.820 ;
        RECT 59.900 214.530 60.150 214.990 ;
        RECT 58.065 214.190 58.625 214.360 ;
        RECT 58.065 214.050 58.235 214.190 ;
        RECT 56.735 213.880 58.235 214.050 ;
        RECT 58.930 214.020 59.390 214.310 ;
        RECT 56.205 213.540 57.895 213.710 ;
        RECT 55.865 213.120 56.220 213.340 ;
        RECT 56.390 212.830 56.560 213.540 ;
        RECT 56.765 213.120 57.555 213.370 ;
        RECT 57.725 213.360 57.895 213.540 ;
        RECT 58.065 213.190 58.235 213.880 ;
        RECT 54.505 212.440 54.835 212.800 ;
        RECT 55.005 212.660 55.500 212.830 ;
        RECT 55.705 212.660 56.560 212.830 ;
        RECT 57.435 212.440 57.765 212.900 ;
        RECT 57.975 212.800 58.235 213.190 ;
        RECT 58.425 214.010 59.390 214.020 ;
        RECT 59.560 214.100 59.730 214.480 ;
        RECT 60.320 214.440 60.490 214.730 ;
        RECT 60.670 214.610 61.000 214.990 ;
        RECT 60.320 214.270 61.120 214.440 ;
        RECT 58.425 213.850 59.100 214.010 ;
        RECT 59.560 213.930 60.780 214.100 ;
        RECT 58.425 213.060 58.635 213.850 ;
        RECT 59.560 213.840 59.730 213.930 ;
        RECT 58.805 213.060 59.155 213.680 ;
        RECT 59.325 213.670 59.730 213.840 ;
        RECT 59.325 212.890 59.495 213.670 ;
        RECT 59.665 213.220 59.885 213.500 ;
        RECT 60.065 213.390 60.605 213.760 ;
        RECT 60.950 213.680 61.120 214.270 ;
        RECT 61.340 213.850 61.645 214.990 ;
        RECT 61.815 213.800 62.070 214.680 ;
        RECT 60.950 213.650 61.690 213.680 ;
        RECT 59.665 213.050 60.195 213.220 ;
        RECT 57.975 212.630 58.325 212.800 ;
        RECT 58.545 212.610 59.495 212.890 ;
        RECT 59.665 212.440 59.855 212.880 ;
        RECT 60.025 212.820 60.195 213.050 ;
        RECT 60.365 212.990 60.605 213.390 ;
        RECT 60.775 213.350 61.690 213.650 ;
        RECT 60.775 213.175 61.100 213.350 ;
        RECT 60.775 212.820 61.095 213.175 ;
        RECT 61.860 213.150 62.070 213.800 ;
        RECT 60.025 212.650 61.095 212.820 ;
        RECT 61.340 212.440 61.645 212.900 ;
        RECT 61.815 212.620 62.070 213.150 ;
        RECT 62.250 213.850 62.585 214.820 ;
        RECT 62.755 213.850 62.925 214.990 ;
        RECT 63.095 214.650 65.125 214.820 ;
        RECT 62.250 213.180 62.420 213.850 ;
        RECT 63.095 213.680 63.265 214.650 ;
        RECT 62.590 213.350 62.845 213.680 ;
        RECT 63.070 213.350 63.265 213.680 ;
        RECT 63.435 214.310 64.560 214.480 ;
        RECT 62.675 213.180 62.845 213.350 ;
        RECT 63.435 213.180 63.605 214.310 ;
        RECT 62.250 212.610 62.505 213.180 ;
        RECT 62.675 213.010 63.605 213.180 ;
        RECT 63.775 213.970 64.785 214.140 ;
        RECT 63.775 213.170 63.945 213.970 ;
        RECT 64.150 213.290 64.425 213.770 ;
        RECT 64.145 213.120 64.425 213.290 ;
        RECT 63.430 212.975 63.605 213.010 ;
        RECT 62.675 212.440 63.005 212.840 ;
        RECT 63.430 212.610 63.960 212.975 ;
        RECT 64.150 212.610 64.425 213.120 ;
        RECT 64.595 212.610 64.785 213.970 ;
        RECT 64.955 213.985 65.125 214.650 ;
        RECT 65.295 214.230 65.465 214.990 ;
        RECT 65.700 214.230 66.215 214.640 ;
        RECT 64.955 213.795 65.705 213.985 ;
        RECT 65.875 213.420 66.215 214.230 ;
        RECT 66.850 214.320 67.105 214.820 ;
        RECT 67.275 214.490 67.605 214.990 ;
        RECT 66.850 214.150 67.600 214.320 ;
        RECT 64.985 213.250 66.215 213.420 ;
        RECT 66.850 213.330 67.200 213.980 ;
        RECT 64.965 212.440 65.475 212.975 ;
        RECT 65.695 212.645 65.940 213.250 ;
        RECT 67.370 213.160 67.600 214.150 ;
        RECT 66.850 212.990 67.600 213.160 ;
        RECT 66.850 212.700 67.105 212.990 ;
        RECT 67.275 212.440 67.605 212.820 ;
        RECT 67.775 212.700 67.945 214.820 ;
        RECT 68.115 214.020 68.440 214.805 ;
        RECT 68.610 214.530 68.860 214.990 ;
        RECT 69.030 214.490 69.280 214.820 ;
        RECT 69.495 214.490 70.175 214.820 ;
        RECT 69.030 214.360 69.200 214.490 ;
        RECT 68.805 214.190 69.200 214.360 ;
        RECT 68.175 212.970 68.635 214.020 ;
        RECT 68.805 212.830 68.975 214.190 ;
        RECT 69.370 213.930 69.835 214.320 ;
        RECT 69.145 213.120 69.495 213.740 ;
        RECT 69.665 213.340 69.835 213.930 ;
        RECT 70.005 213.710 70.175 214.490 ;
        RECT 70.345 214.390 70.515 214.730 ;
        RECT 70.750 214.560 71.080 214.990 ;
        RECT 71.250 214.390 71.420 214.730 ;
        RECT 71.715 214.530 72.085 214.990 ;
        RECT 70.345 214.220 71.420 214.390 ;
        RECT 72.255 214.360 72.425 214.820 ;
        RECT 72.660 214.480 73.530 214.820 ;
        RECT 73.700 214.530 73.950 214.990 ;
        RECT 71.865 214.190 72.425 214.360 ;
        RECT 71.865 214.050 72.035 214.190 ;
        RECT 70.535 213.880 72.035 214.050 ;
        RECT 72.730 214.020 73.190 214.310 ;
        RECT 70.005 213.540 71.695 213.710 ;
        RECT 69.665 213.120 70.020 213.340 ;
        RECT 70.190 212.830 70.360 213.540 ;
        RECT 70.565 213.120 71.355 213.370 ;
        RECT 71.525 213.360 71.695 213.540 ;
        RECT 71.865 213.190 72.035 213.880 ;
        RECT 68.305 212.440 68.635 212.800 ;
        RECT 68.805 212.660 69.300 212.830 ;
        RECT 69.505 212.660 70.360 212.830 ;
        RECT 71.235 212.440 71.565 212.900 ;
        RECT 71.775 212.800 72.035 213.190 ;
        RECT 72.225 214.010 73.190 214.020 ;
        RECT 73.360 214.100 73.530 214.480 ;
        RECT 74.120 214.440 74.290 214.730 ;
        RECT 74.470 214.610 74.800 214.990 ;
        RECT 74.120 214.270 74.920 214.440 ;
        RECT 72.225 213.850 72.900 214.010 ;
        RECT 73.360 213.930 74.580 214.100 ;
        RECT 72.225 213.060 72.435 213.850 ;
        RECT 73.360 213.840 73.530 213.930 ;
        RECT 72.605 213.060 72.955 213.680 ;
        RECT 73.125 213.670 73.530 213.840 ;
        RECT 73.125 212.890 73.295 213.670 ;
        RECT 73.465 213.220 73.685 213.500 ;
        RECT 73.865 213.390 74.405 213.760 ;
        RECT 74.750 213.680 74.920 214.270 ;
        RECT 75.140 213.850 75.445 214.990 ;
        RECT 75.615 213.800 75.865 214.680 ;
        RECT 76.035 213.850 76.285 214.990 ;
        RECT 76.545 213.850 76.775 214.990 ;
        RECT 76.945 213.840 77.275 214.820 ;
        RECT 77.445 213.850 77.655 214.990 ;
        RECT 74.750 213.650 75.490 213.680 ;
        RECT 73.465 213.050 73.995 213.220 ;
        RECT 71.775 212.630 72.125 212.800 ;
        RECT 72.345 212.610 73.295 212.890 ;
        RECT 73.465 212.440 73.655 212.880 ;
        RECT 73.825 212.820 73.995 213.050 ;
        RECT 74.165 212.990 74.405 213.390 ;
        RECT 74.575 213.350 75.490 213.650 ;
        RECT 74.575 213.175 74.900 213.350 ;
        RECT 74.575 212.820 74.895 213.175 ;
        RECT 75.660 213.150 75.865 213.800 ;
        RECT 76.525 213.430 76.855 213.680 ;
        RECT 73.825 212.650 74.895 212.820 ;
        RECT 75.140 212.440 75.445 212.900 ;
        RECT 75.615 212.620 75.865 213.150 ;
        RECT 76.035 212.440 76.285 213.195 ;
        RECT 76.545 212.440 76.775 213.260 ;
        RECT 77.025 213.240 77.275 213.840 ;
        RECT 78.345 213.825 78.635 214.990 ;
        RECT 78.855 213.850 79.105 214.990 ;
        RECT 79.275 213.800 79.525 214.680 ;
        RECT 79.695 213.850 80.000 214.990 ;
        RECT 80.340 214.610 80.670 214.990 ;
        RECT 80.850 214.440 81.020 214.730 ;
        RECT 81.190 214.530 81.440 214.990 ;
        RECT 80.220 214.270 81.020 214.440 ;
        RECT 81.610 214.480 82.480 214.820 ;
        RECT 76.945 212.610 77.275 213.240 ;
        RECT 77.445 212.440 77.655 213.260 ;
        RECT 78.345 212.440 78.635 213.165 ;
        RECT 78.855 212.440 79.105 213.195 ;
        RECT 79.275 213.150 79.480 213.800 ;
        RECT 80.220 213.680 80.390 214.270 ;
        RECT 81.610 214.100 81.780 214.480 ;
        RECT 82.715 214.360 82.885 214.820 ;
        RECT 83.055 214.530 83.425 214.990 ;
        RECT 83.720 214.390 83.890 214.730 ;
        RECT 84.060 214.560 84.390 214.990 ;
        RECT 84.625 214.390 84.795 214.730 ;
        RECT 80.560 213.930 81.780 214.100 ;
        RECT 81.950 214.020 82.410 214.310 ;
        RECT 82.715 214.190 83.275 214.360 ;
        RECT 83.720 214.220 84.795 214.390 ;
        RECT 84.965 214.490 85.645 214.820 ;
        RECT 85.860 214.490 86.110 214.820 ;
        RECT 86.280 214.530 86.530 214.990 ;
        RECT 83.105 214.050 83.275 214.190 ;
        RECT 81.950 214.010 82.915 214.020 ;
        RECT 81.610 213.840 81.780 213.930 ;
        RECT 82.240 213.850 82.915 214.010 ;
        RECT 79.650 213.650 80.390 213.680 ;
        RECT 79.650 213.350 80.565 213.650 ;
        RECT 80.240 213.175 80.565 213.350 ;
        RECT 79.275 212.620 79.525 213.150 ;
        RECT 79.695 212.440 80.000 212.900 ;
        RECT 80.245 212.820 80.565 213.175 ;
        RECT 80.735 213.390 81.275 213.760 ;
        RECT 81.610 213.670 82.015 213.840 ;
        RECT 80.735 212.990 80.975 213.390 ;
        RECT 81.455 213.220 81.675 213.500 ;
        RECT 81.145 213.050 81.675 213.220 ;
        RECT 81.145 212.820 81.315 213.050 ;
        RECT 81.845 212.890 82.015 213.670 ;
        RECT 82.185 213.060 82.535 213.680 ;
        RECT 82.705 213.060 82.915 213.850 ;
        RECT 83.105 213.880 84.605 214.050 ;
        RECT 83.105 213.190 83.275 213.880 ;
        RECT 84.965 213.710 85.135 214.490 ;
        RECT 85.940 214.360 86.110 214.490 ;
        RECT 83.445 213.540 85.135 213.710 ;
        RECT 85.305 213.930 85.770 214.320 ;
        RECT 85.940 214.190 86.335 214.360 ;
        RECT 83.445 213.360 83.615 213.540 ;
        RECT 80.245 212.650 81.315 212.820 ;
        RECT 81.485 212.440 81.675 212.880 ;
        RECT 81.845 212.610 82.795 212.890 ;
        RECT 83.105 212.800 83.365 213.190 ;
        RECT 83.785 213.120 84.575 213.370 ;
        RECT 83.015 212.630 83.365 212.800 ;
        RECT 83.575 212.440 83.905 212.900 ;
        RECT 84.780 212.830 84.950 213.540 ;
        RECT 85.305 213.340 85.475 213.930 ;
        RECT 85.120 213.120 85.475 213.340 ;
        RECT 85.645 213.120 85.995 213.740 ;
        RECT 86.165 212.830 86.335 214.190 ;
        RECT 86.700 214.020 87.025 214.805 ;
        RECT 86.505 212.970 86.965 214.020 ;
        RECT 84.780 212.660 85.635 212.830 ;
        RECT 85.840 212.660 86.335 212.830 ;
        RECT 86.505 212.440 86.835 212.800 ;
        RECT 87.195 212.700 87.365 214.820 ;
        RECT 87.535 214.490 87.865 214.990 ;
        RECT 88.035 214.320 88.290 214.820 ;
        RECT 87.540 214.150 88.290 214.320 ;
        RECT 88.470 214.320 88.725 214.820 ;
        RECT 88.895 214.490 89.225 214.990 ;
        RECT 88.470 214.150 89.220 214.320 ;
        RECT 87.540 213.160 87.770 214.150 ;
        RECT 87.940 213.330 88.290 213.980 ;
        RECT 88.470 213.330 88.820 213.980 ;
        RECT 88.990 213.160 89.220 214.150 ;
        RECT 87.540 212.990 88.290 213.160 ;
        RECT 87.535 212.440 87.865 212.820 ;
        RECT 88.035 212.700 88.290 212.990 ;
        RECT 88.470 212.990 89.220 213.160 ;
        RECT 88.470 212.700 88.725 212.990 ;
        RECT 88.895 212.440 89.225 212.820 ;
        RECT 89.395 212.700 89.565 214.820 ;
        RECT 89.735 214.020 90.060 214.805 ;
        RECT 90.230 214.530 90.480 214.990 ;
        RECT 90.650 214.490 90.900 214.820 ;
        RECT 91.115 214.490 91.795 214.820 ;
        RECT 90.650 214.360 90.820 214.490 ;
        RECT 90.425 214.190 90.820 214.360 ;
        RECT 89.795 212.970 90.255 214.020 ;
        RECT 90.425 212.830 90.595 214.190 ;
        RECT 90.990 213.930 91.455 214.320 ;
        RECT 90.765 213.120 91.115 213.740 ;
        RECT 91.285 213.340 91.455 213.930 ;
        RECT 91.625 213.710 91.795 214.490 ;
        RECT 91.965 214.390 92.135 214.730 ;
        RECT 92.370 214.560 92.700 214.990 ;
        RECT 92.870 214.390 93.040 214.730 ;
        RECT 93.335 214.530 93.705 214.990 ;
        RECT 91.965 214.220 93.040 214.390 ;
        RECT 93.875 214.360 94.045 214.820 ;
        RECT 94.280 214.480 95.150 214.820 ;
        RECT 95.320 214.530 95.570 214.990 ;
        RECT 93.485 214.190 94.045 214.360 ;
        RECT 93.485 214.050 93.655 214.190 ;
        RECT 92.155 213.880 93.655 214.050 ;
        RECT 94.350 214.020 94.810 214.310 ;
        RECT 91.625 213.540 93.315 213.710 ;
        RECT 91.285 213.120 91.640 213.340 ;
        RECT 91.810 212.830 91.980 213.540 ;
        RECT 92.185 213.120 92.975 213.370 ;
        RECT 93.145 213.360 93.315 213.540 ;
        RECT 93.485 213.190 93.655 213.880 ;
        RECT 89.925 212.440 90.255 212.800 ;
        RECT 90.425 212.660 90.920 212.830 ;
        RECT 91.125 212.660 91.980 212.830 ;
        RECT 92.855 212.440 93.185 212.900 ;
        RECT 93.395 212.800 93.655 213.190 ;
        RECT 93.845 214.010 94.810 214.020 ;
        RECT 94.980 214.100 95.150 214.480 ;
        RECT 95.740 214.440 95.910 214.730 ;
        RECT 96.090 214.610 96.420 214.990 ;
        RECT 95.740 214.270 96.540 214.440 ;
        RECT 93.845 213.850 94.520 214.010 ;
        RECT 94.980 213.930 96.200 214.100 ;
        RECT 93.845 213.060 94.055 213.850 ;
        RECT 94.980 213.840 95.150 213.930 ;
        RECT 94.225 213.060 94.575 213.680 ;
        RECT 94.745 213.670 95.150 213.840 ;
        RECT 94.745 212.890 94.915 213.670 ;
        RECT 95.085 213.220 95.305 213.500 ;
        RECT 95.485 213.390 96.025 213.760 ;
        RECT 96.370 213.680 96.540 214.270 ;
        RECT 96.760 213.850 97.065 214.990 ;
        RECT 97.235 213.800 97.490 214.680 ;
        RECT 97.865 214.320 98.145 214.990 ;
        RECT 98.315 214.100 98.615 214.650 ;
        RECT 98.815 214.270 99.145 214.990 ;
        RECT 99.335 214.270 99.795 214.820 ;
        RECT 96.370 213.650 97.110 213.680 ;
        RECT 95.085 213.050 95.615 213.220 ;
        RECT 93.395 212.630 93.745 212.800 ;
        RECT 93.965 212.610 94.915 212.890 ;
        RECT 95.085 212.440 95.275 212.880 ;
        RECT 95.445 212.820 95.615 213.050 ;
        RECT 95.785 212.990 96.025 213.390 ;
        RECT 96.195 213.350 97.110 213.650 ;
        RECT 96.195 213.175 96.520 213.350 ;
        RECT 96.195 212.820 96.515 213.175 ;
        RECT 97.280 213.150 97.490 213.800 ;
        RECT 97.680 213.680 97.945 214.040 ;
        RECT 98.315 213.930 99.255 214.100 ;
        RECT 99.085 213.680 99.255 213.930 ;
        RECT 97.680 213.430 98.355 213.680 ;
        RECT 98.575 213.430 98.915 213.680 ;
        RECT 99.085 213.350 99.375 213.680 ;
        RECT 99.085 213.260 99.255 213.350 ;
        RECT 95.445 212.650 96.515 212.820 ;
        RECT 96.760 212.440 97.065 212.900 ;
        RECT 97.235 212.620 97.490 213.150 ;
        RECT 97.865 213.070 99.255 213.260 ;
        RECT 97.865 212.710 98.195 213.070 ;
        RECT 99.545 212.900 99.795 214.270 ;
        RECT 98.815 212.440 99.065 212.900 ;
        RECT 99.235 212.610 99.795 212.900 ;
        RECT 99.970 213.850 100.305 214.820 ;
        RECT 100.475 213.850 100.645 214.990 ;
        RECT 100.815 214.650 102.845 214.820 ;
        RECT 99.970 213.180 100.140 213.850 ;
        RECT 100.815 213.680 100.985 214.650 ;
        RECT 100.310 213.350 100.565 213.680 ;
        RECT 100.790 213.350 100.985 213.680 ;
        RECT 101.155 214.310 102.280 214.480 ;
        RECT 100.395 213.180 100.565 213.350 ;
        RECT 101.155 213.180 101.325 214.310 ;
        RECT 99.970 212.610 100.225 213.180 ;
        RECT 100.395 213.010 101.325 213.180 ;
        RECT 101.495 213.970 102.505 214.140 ;
        RECT 101.495 213.170 101.665 213.970 ;
        RECT 101.870 213.630 102.145 213.770 ;
        RECT 101.865 213.460 102.145 213.630 ;
        RECT 101.150 212.975 101.325 213.010 ;
        RECT 100.395 212.440 100.725 212.840 ;
        RECT 101.150 212.610 101.680 212.975 ;
        RECT 101.870 212.610 102.145 213.460 ;
        RECT 102.315 212.610 102.505 213.970 ;
        RECT 102.675 213.985 102.845 214.650 ;
        RECT 103.015 214.230 103.185 214.990 ;
        RECT 103.420 214.230 103.935 214.640 ;
        RECT 102.675 213.795 103.425 213.985 ;
        RECT 103.595 213.420 103.935 214.230 ;
        RECT 104.105 213.825 104.395 214.990 ;
        RECT 102.705 213.250 103.935 213.420 ;
        RECT 102.685 212.440 103.195 212.975 ;
        RECT 103.415 212.645 103.660 213.250 ;
        RECT 104.105 212.440 104.395 213.165 ;
        RECT 104.575 212.620 104.835 214.810 ;
        RECT 105.005 214.260 105.345 214.990 ;
        RECT 105.525 214.080 105.795 214.810 ;
        RECT 105.025 213.860 105.795 214.080 ;
        RECT 105.975 214.100 106.205 214.810 ;
        RECT 106.375 214.280 106.705 214.990 ;
        RECT 106.875 214.100 107.135 214.810 ;
        RECT 107.330 214.565 107.665 214.990 ;
        RECT 107.835 214.385 108.020 214.790 ;
        RECT 105.975 213.860 107.135 214.100 ;
        RECT 107.355 214.210 108.020 214.385 ;
        RECT 108.225 214.210 108.555 214.990 ;
        RECT 105.025 213.190 105.315 213.860 ;
        RECT 105.495 213.370 105.960 213.680 ;
        RECT 106.140 213.370 106.665 213.680 ;
        RECT 105.025 212.990 106.255 213.190 ;
        RECT 105.095 212.440 105.765 212.810 ;
        RECT 105.945 212.620 106.255 212.990 ;
        RECT 106.435 212.730 106.665 213.370 ;
        RECT 106.845 213.350 107.145 213.680 ;
        RECT 107.355 213.180 107.695 214.210 ;
        RECT 108.725 214.020 108.995 214.790 ;
        RECT 107.865 213.850 108.995 214.020 ;
        RECT 109.165 213.900 110.835 214.990 ;
        RECT 107.865 213.350 108.115 213.850 ;
        RECT 106.845 212.440 107.135 213.170 ;
        RECT 107.355 213.010 108.040 213.180 ;
        RECT 108.295 213.100 108.655 213.680 ;
        RECT 107.330 212.440 107.665 212.840 ;
        RECT 107.835 212.610 108.040 213.010 ;
        RECT 108.825 212.940 108.995 213.850 ;
        RECT 108.250 212.440 108.525 212.920 ;
        RECT 108.735 212.610 108.995 212.940 ;
        RECT 109.165 213.210 109.915 213.730 ;
        RECT 110.085 213.380 110.835 213.900 ;
        RECT 111.010 213.850 111.345 214.820 ;
        RECT 111.515 213.850 111.685 214.990 ;
        RECT 111.855 214.650 113.885 214.820 ;
        RECT 109.165 212.440 110.835 213.210 ;
        RECT 111.010 213.180 111.180 213.850 ;
        RECT 111.855 213.680 112.025 214.650 ;
        RECT 111.350 213.350 111.605 213.680 ;
        RECT 111.830 213.350 112.025 213.680 ;
        RECT 112.195 214.310 113.320 214.480 ;
        RECT 111.435 213.180 111.605 213.350 ;
        RECT 112.195 213.180 112.365 214.310 ;
        RECT 111.010 212.610 111.265 213.180 ;
        RECT 111.435 213.010 112.365 213.180 ;
        RECT 112.535 213.970 113.545 214.140 ;
        RECT 112.535 213.170 112.705 213.970 ;
        RECT 112.190 212.975 112.365 213.010 ;
        RECT 111.435 212.440 111.765 212.840 ;
        RECT 112.190 212.610 112.720 212.975 ;
        RECT 112.910 212.950 113.185 213.770 ;
        RECT 112.905 212.780 113.185 212.950 ;
        RECT 112.910 212.610 113.185 212.780 ;
        RECT 113.355 212.610 113.545 213.970 ;
        RECT 113.715 213.985 113.885 214.650 ;
        RECT 114.055 214.230 114.225 214.990 ;
        RECT 114.460 214.230 114.975 214.640 ;
        RECT 113.715 213.795 114.465 213.985 ;
        RECT 114.635 213.420 114.975 214.230 ;
        RECT 116.105 213.850 116.335 214.990 ;
        RECT 116.505 213.840 116.835 214.820 ;
        RECT 117.005 213.850 117.215 214.990 ;
        RECT 117.445 214.150 117.875 214.990 ;
        RECT 118.465 214.490 118.715 214.990 ;
        RECT 118.985 214.650 120.110 214.820 ;
        RECT 118.985 214.490 119.235 214.650 ;
        RECT 119.785 214.480 120.110 214.650 ;
        RECT 120.280 214.490 120.530 214.990 ;
        RECT 120.700 214.480 120.950 214.820 ;
        RECT 118.045 214.320 118.295 214.480 ;
        RECT 119.405 214.320 119.615 214.480 ;
        RECT 118.045 214.150 119.615 214.320 ;
        RECT 121.260 214.320 121.510 214.820 ;
        RECT 121.680 214.490 121.930 214.990 ;
        RECT 122.100 214.320 122.350 214.820 ;
        RECT 122.520 214.490 122.770 214.990 ;
        RECT 122.940 214.320 123.255 214.820 ;
        RECT 123.925 214.530 124.140 214.990 ;
        RECT 124.310 214.360 124.640 214.820 ;
        RECT 121.260 214.310 123.255 214.320 ;
        RECT 118.045 213.980 118.295 214.150 ;
        RECT 119.860 214.140 123.255 214.310 ;
        RECT 119.860 213.980 120.030 214.140 ;
        RECT 116.085 213.430 116.415 213.680 ;
        RECT 113.745 213.250 114.975 213.420 ;
        RECT 113.725 212.440 114.235 212.975 ;
        RECT 114.455 212.645 114.700 213.250 ;
        RECT 116.105 212.440 116.335 213.260 ;
        RECT 116.585 213.240 116.835 213.840 ;
        RECT 117.445 213.770 118.295 213.980 ;
        RECT 118.535 213.810 120.030 213.980 ;
        RECT 116.505 212.610 116.835 213.240 ;
        RECT 117.005 212.440 117.215 213.260 ;
        RECT 117.445 212.830 117.835 213.770 ;
        RECT 118.535 213.600 118.705 213.810 ;
        RECT 120.240 213.800 122.550 213.970 ;
        RECT 120.240 213.640 120.410 213.800 ;
        RECT 118.045 213.430 118.705 213.600 ;
        RECT 119.385 213.430 120.410 213.640 ;
        RECT 122.380 213.640 122.550 213.800 ;
        RECT 120.635 213.430 122.085 213.630 ;
        RECT 122.380 213.430 122.855 213.640 ;
        RECT 118.005 213.080 120.570 213.260 ;
        RECT 118.005 213.000 118.335 213.080 ;
        RECT 117.445 212.660 118.755 212.830 ;
        RECT 119.025 212.440 119.195 212.910 ;
        RECT 119.365 212.610 119.730 213.080 ;
        RECT 119.900 212.440 120.070 212.910 ;
        RECT 120.240 212.610 120.570 213.080 ;
        RECT 120.740 212.440 120.910 213.260 ;
        RECT 121.220 213.080 122.310 213.260 ;
        RECT 123.025 213.250 123.255 214.140 ;
        RECT 121.220 212.610 121.550 213.080 ;
        RECT 121.720 212.440 121.890 212.910 ;
        RECT 122.060 212.830 122.310 213.080 ;
        RECT 122.480 213.000 123.255 213.250 ;
        RECT 123.470 214.190 124.640 214.360 ;
        RECT 124.810 214.190 125.060 214.990 ;
        RECT 123.470 212.900 123.840 214.190 ;
        RECT 125.270 214.020 125.550 214.180 ;
        RECT 124.215 213.850 125.550 214.020 ;
        RECT 124.215 213.680 124.385 213.850 ;
        RECT 124.010 213.430 124.385 213.680 ;
        RECT 124.555 213.430 125.030 213.670 ;
        RECT 125.200 213.430 125.550 213.670 ;
        RECT 124.215 213.260 124.385 213.430 ;
        RECT 124.215 213.090 125.550 213.260 ;
        RECT 122.060 212.610 123.235 212.830 ;
        RECT 123.470 212.610 124.220 212.900 ;
        RECT 124.730 212.440 125.060 212.900 ;
        RECT 125.280 212.880 125.550 213.090 ;
        RECT 126.195 212.620 126.455 214.810 ;
        RECT 126.625 214.260 126.965 214.990 ;
        RECT 127.145 214.080 127.415 214.810 ;
        RECT 126.645 213.860 127.415 214.080 ;
        RECT 127.595 214.100 127.825 214.810 ;
        RECT 127.995 214.280 128.325 214.990 ;
        RECT 128.495 214.100 128.755 214.810 ;
        RECT 127.595 213.860 128.755 214.100 ;
        RECT 126.645 213.190 126.935 213.860 ;
        RECT 129.865 213.825 130.155 214.990 ;
        RECT 130.330 214.320 130.585 214.820 ;
        RECT 130.755 214.490 131.085 214.990 ;
        RECT 130.330 214.150 131.080 214.320 ;
        RECT 127.115 213.370 127.580 213.680 ;
        RECT 127.760 213.370 128.285 213.680 ;
        RECT 126.645 212.990 127.875 213.190 ;
        RECT 126.715 212.440 127.385 212.810 ;
        RECT 127.565 212.620 127.875 212.990 ;
        RECT 128.055 212.730 128.285 213.370 ;
        RECT 128.465 213.350 128.765 213.680 ;
        RECT 130.330 213.330 130.680 213.980 ;
        RECT 128.465 212.440 128.755 213.170 ;
        RECT 129.865 212.440 130.155 213.165 ;
        RECT 130.850 213.160 131.080 214.150 ;
        RECT 130.330 212.990 131.080 213.160 ;
        RECT 130.330 212.700 130.585 212.990 ;
        RECT 130.755 212.440 131.085 212.820 ;
        RECT 131.255 212.700 131.425 214.820 ;
        RECT 131.595 214.020 131.920 214.805 ;
        RECT 132.090 214.530 132.340 214.990 ;
        RECT 132.510 214.490 132.760 214.820 ;
        RECT 132.975 214.490 133.655 214.820 ;
        RECT 132.510 214.360 132.680 214.490 ;
        RECT 132.285 214.190 132.680 214.360 ;
        RECT 131.655 212.970 132.115 214.020 ;
        RECT 132.285 212.830 132.455 214.190 ;
        RECT 132.850 213.930 133.315 214.320 ;
        RECT 132.625 213.120 132.975 213.740 ;
        RECT 133.145 213.340 133.315 213.930 ;
        RECT 133.485 213.710 133.655 214.490 ;
        RECT 133.825 214.390 133.995 214.730 ;
        RECT 134.230 214.560 134.560 214.990 ;
        RECT 134.730 214.390 134.900 214.730 ;
        RECT 135.195 214.530 135.565 214.990 ;
        RECT 133.825 214.220 134.900 214.390 ;
        RECT 135.735 214.360 135.905 214.820 ;
        RECT 136.140 214.480 137.010 214.820 ;
        RECT 137.180 214.530 137.430 214.990 ;
        RECT 135.345 214.190 135.905 214.360 ;
        RECT 135.345 214.050 135.515 214.190 ;
        RECT 134.015 213.880 135.515 214.050 ;
        RECT 136.210 214.020 136.670 214.310 ;
        RECT 133.485 213.540 135.175 213.710 ;
        RECT 133.145 213.120 133.500 213.340 ;
        RECT 133.670 212.830 133.840 213.540 ;
        RECT 134.045 213.120 134.835 213.370 ;
        RECT 135.005 213.360 135.175 213.540 ;
        RECT 135.345 213.190 135.515 213.880 ;
        RECT 131.785 212.440 132.115 212.800 ;
        RECT 132.285 212.660 132.780 212.830 ;
        RECT 132.985 212.660 133.840 212.830 ;
        RECT 134.715 212.440 135.045 212.900 ;
        RECT 135.255 212.800 135.515 213.190 ;
        RECT 135.705 214.010 136.670 214.020 ;
        RECT 136.840 214.100 137.010 214.480 ;
        RECT 137.600 214.440 137.770 214.730 ;
        RECT 137.950 214.610 138.280 214.990 ;
        RECT 137.600 214.270 138.400 214.440 ;
        RECT 135.705 213.850 136.380 214.010 ;
        RECT 136.840 213.930 138.060 214.100 ;
        RECT 135.705 213.060 135.915 213.850 ;
        RECT 136.840 213.840 137.010 213.930 ;
        RECT 136.085 213.060 136.435 213.680 ;
        RECT 136.605 213.670 137.010 213.840 ;
        RECT 136.605 212.890 136.775 213.670 ;
        RECT 136.945 213.220 137.165 213.500 ;
        RECT 137.345 213.390 137.885 213.760 ;
        RECT 138.230 213.680 138.400 214.270 ;
        RECT 138.620 213.850 138.925 214.990 ;
        RECT 139.095 213.800 139.350 214.680 ;
        RECT 139.530 213.840 139.790 214.990 ;
        RECT 139.965 213.915 140.220 214.820 ;
        RECT 140.390 214.230 140.720 214.990 ;
        RECT 140.935 214.060 141.105 214.820 ;
        RECT 138.230 213.650 138.970 213.680 ;
        RECT 136.945 213.050 137.475 213.220 ;
        RECT 135.255 212.630 135.605 212.800 ;
        RECT 135.825 212.610 136.775 212.890 ;
        RECT 136.945 212.440 137.135 212.880 ;
        RECT 137.305 212.820 137.475 213.050 ;
        RECT 137.645 212.990 137.885 213.390 ;
        RECT 138.055 213.350 138.970 213.650 ;
        RECT 138.055 213.175 138.380 213.350 ;
        RECT 138.055 212.820 138.375 213.175 ;
        RECT 139.140 213.150 139.350 213.800 ;
        RECT 137.305 212.650 138.375 212.820 ;
        RECT 138.620 212.440 138.925 212.900 ;
        RECT 139.095 212.620 139.350 213.150 ;
        RECT 139.530 212.440 139.790 213.280 ;
        RECT 139.965 213.185 140.135 213.915 ;
        RECT 140.390 213.890 141.105 214.060 ;
        RECT 141.365 213.915 141.635 214.820 ;
        RECT 141.805 214.230 142.135 214.990 ;
        RECT 142.315 214.060 142.495 214.820 ;
        RECT 140.390 213.680 140.560 213.890 ;
        RECT 140.305 213.350 140.560 213.680 ;
        RECT 139.965 212.610 140.220 213.185 ;
        RECT 140.390 213.160 140.560 213.350 ;
        RECT 140.840 213.340 141.195 213.710 ;
        RECT 140.390 212.990 141.105 213.160 ;
        RECT 140.390 212.440 140.720 212.820 ;
        RECT 140.935 212.610 141.105 212.990 ;
        RECT 141.365 213.115 141.545 213.915 ;
        RECT 141.820 213.890 142.495 214.060 ;
        RECT 142.835 214.060 143.005 214.820 ;
        RECT 143.220 214.230 143.550 214.990 ;
        RECT 142.835 213.890 143.550 214.060 ;
        RECT 143.720 213.915 143.975 214.820 ;
        RECT 141.820 213.745 141.990 213.890 ;
        RECT 141.715 213.415 141.990 213.745 ;
        RECT 141.820 213.160 141.990 213.415 ;
        RECT 142.215 213.340 142.555 213.710 ;
        RECT 142.745 213.340 143.100 213.710 ;
        RECT 143.380 213.680 143.550 213.890 ;
        RECT 143.380 213.350 143.635 213.680 ;
        RECT 143.380 213.160 143.550 213.350 ;
        RECT 143.805 213.185 143.975 213.915 ;
        RECT 144.150 213.840 144.410 214.990 ;
        RECT 144.675 214.060 144.845 214.820 ;
        RECT 145.060 214.230 145.390 214.990 ;
        RECT 144.675 213.890 145.390 214.060 ;
        RECT 145.560 213.915 145.815 214.820 ;
        RECT 144.585 213.340 144.940 213.710 ;
        RECT 145.220 213.680 145.390 213.890 ;
        RECT 145.220 213.350 145.475 213.680 ;
        RECT 141.365 212.610 141.625 213.115 ;
        RECT 141.820 212.990 142.485 213.160 ;
        RECT 141.805 212.440 142.135 212.820 ;
        RECT 142.315 212.610 142.485 212.990 ;
        RECT 142.835 212.990 143.550 213.160 ;
        RECT 142.835 212.610 143.005 212.990 ;
        RECT 143.220 212.440 143.550 212.820 ;
        RECT 143.720 212.610 143.975 213.185 ;
        RECT 144.150 212.440 144.410 213.280 ;
        RECT 145.220 213.160 145.390 213.350 ;
        RECT 145.645 213.185 145.815 213.915 ;
        RECT 145.990 213.840 146.250 214.990 ;
        RECT 146.425 213.900 147.635 214.990 ;
        RECT 146.425 213.360 146.945 213.900 ;
        RECT 144.675 212.990 145.390 213.160 ;
        RECT 144.675 212.610 144.845 212.990 ;
        RECT 145.060 212.440 145.390 212.820 ;
        RECT 145.560 212.610 145.815 213.185 ;
        RECT 145.990 212.440 146.250 213.280 ;
        RECT 147.115 213.190 147.635 213.730 ;
        RECT 146.425 212.440 147.635 213.190 ;
        RECT 13.860 212.270 147.720 212.440 ;
        RECT 13.945 211.520 15.155 212.270 ;
        RECT 13.945 210.980 14.465 211.520 ;
        RECT 15.330 211.430 15.590 212.270 ;
        RECT 15.765 211.525 16.020 212.100 ;
        RECT 16.190 211.890 16.520 212.270 ;
        RECT 16.735 211.720 16.905 212.100 ;
        RECT 16.190 211.550 16.905 211.720 ;
        RECT 14.635 210.810 15.155 211.350 ;
        RECT 13.945 209.720 15.155 210.810 ;
        RECT 15.330 209.720 15.590 210.870 ;
        RECT 15.765 210.795 15.935 211.525 ;
        RECT 16.190 211.360 16.360 211.550 ;
        RECT 17.170 211.430 17.430 212.270 ;
        RECT 17.605 211.525 17.860 212.100 ;
        RECT 18.030 211.890 18.360 212.270 ;
        RECT 18.575 211.720 18.745 212.100 ;
        RECT 18.030 211.550 18.745 211.720 ;
        RECT 19.010 211.720 19.265 212.010 ;
        RECT 19.435 211.890 19.765 212.270 ;
        RECT 19.010 211.550 19.760 211.720 ;
        RECT 16.105 211.030 16.360 211.360 ;
        RECT 16.190 210.820 16.360 211.030 ;
        RECT 16.640 211.000 16.995 211.370 ;
        RECT 15.765 209.890 16.020 210.795 ;
        RECT 16.190 210.650 16.905 210.820 ;
        RECT 16.190 209.720 16.520 210.480 ;
        RECT 16.735 209.890 16.905 210.650 ;
        RECT 17.170 209.720 17.430 210.870 ;
        RECT 17.605 210.795 17.775 211.525 ;
        RECT 18.030 211.360 18.200 211.550 ;
        RECT 17.945 211.030 18.200 211.360 ;
        RECT 18.030 210.820 18.200 211.030 ;
        RECT 18.480 211.000 18.835 211.370 ;
        RECT 17.605 209.890 17.860 210.795 ;
        RECT 18.030 210.650 18.745 210.820 ;
        RECT 19.010 210.730 19.360 211.380 ;
        RECT 18.030 209.720 18.360 210.480 ;
        RECT 18.575 209.890 18.745 210.650 ;
        RECT 19.530 210.560 19.760 211.550 ;
        RECT 19.010 210.390 19.760 210.560 ;
        RECT 19.010 209.890 19.265 210.390 ;
        RECT 19.435 209.720 19.765 210.220 ;
        RECT 19.935 209.890 20.105 212.010 ;
        RECT 20.465 211.910 20.795 212.270 ;
        RECT 20.965 211.880 21.460 212.050 ;
        RECT 21.665 211.880 22.520 212.050 ;
        RECT 20.335 210.690 20.795 211.740 ;
        RECT 20.275 209.905 20.600 210.690 ;
        RECT 20.965 210.520 21.135 211.880 ;
        RECT 21.305 210.970 21.655 211.590 ;
        RECT 21.825 211.370 22.180 211.590 ;
        RECT 21.825 210.780 21.995 211.370 ;
        RECT 22.350 211.170 22.520 211.880 ;
        RECT 23.395 211.810 23.725 212.270 ;
        RECT 23.935 211.910 24.285 212.080 ;
        RECT 22.725 211.340 23.515 211.590 ;
        RECT 23.935 211.520 24.195 211.910 ;
        RECT 24.505 211.820 25.455 212.100 ;
        RECT 25.625 211.830 25.815 212.270 ;
        RECT 25.985 211.890 27.055 212.060 ;
        RECT 23.685 211.170 23.855 211.350 ;
        RECT 20.965 210.350 21.360 210.520 ;
        RECT 21.530 210.390 21.995 210.780 ;
        RECT 22.165 211.000 23.855 211.170 ;
        RECT 21.190 210.220 21.360 210.350 ;
        RECT 22.165 210.220 22.335 211.000 ;
        RECT 24.025 210.830 24.195 211.520 ;
        RECT 22.695 210.660 24.195 210.830 ;
        RECT 24.385 210.860 24.595 211.650 ;
        RECT 24.765 211.030 25.115 211.650 ;
        RECT 25.285 211.040 25.455 211.820 ;
        RECT 25.985 211.660 26.155 211.890 ;
        RECT 25.625 211.490 26.155 211.660 ;
        RECT 25.625 211.210 25.845 211.490 ;
        RECT 26.325 211.320 26.565 211.720 ;
        RECT 25.285 210.870 25.690 211.040 ;
        RECT 26.025 210.950 26.565 211.320 ;
        RECT 26.735 211.535 27.055 211.890 ;
        RECT 26.735 211.280 27.060 211.535 ;
        RECT 27.255 211.460 27.425 212.270 ;
        RECT 27.595 211.620 27.925 212.100 ;
        RECT 28.095 211.800 28.265 212.270 ;
        RECT 28.435 211.620 28.765 212.100 ;
        RECT 28.935 211.800 29.105 212.270 ;
        RECT 27.595 211.450 29.360 211.620 ;
        RECT 26.735 211.070 28.765 211.280 ;
        RECT 26.735 211.060 27.080 211.070 ;
        RECT 24.385 210.700 25.060 210.860 ;
        RECT 25.520 210.780 25.690 210.870 ;
        RECT 24.385 210.690 25.350 210.700 ;
        RECT 24.025 210.520 24.195 210.660 ;
        RECT 20.770 209.720 21.020 210.180 ;
        RECT 21.190 209.890 21.440 210.220 ;
        RECT 21.655 209.890 22.335 210.220 ;
        RECT 22.505 210.320 23.580 210.490 ;
        RECT 24.025 210.350 24.585 210.520 ;
        RECT 24.890 210.400 25.350 210.690 ;
        RECT 25.520 210.610 26.740 210.780 ;
        RECT 22.505 209.980 22.675 210.320 ;
        RECT 22.910 209.720 23.240 210.150 ;
        RECT 23.410 209.980 23.580 210.320 ;
        RECT 23.875 209.720 24.245 210.180 ;
        RECT 24.415 209.890 24.585 210.350 ;
        RECT 25.520 210.230 25.690 210.610 ;
        RECT 26.910 210.440 27.080 211.060 ;
        RECT 28.950 210.900 29.360 211.450 ;
        RECT 29.585 211.500 31.255 212.270 ;
        RECT 31.430 211.530 31.685 212.100 ;
        RECT 31.855 211.870 32.185 212.270 ;
        RECT 32.610 211.735 33.140 212.100 ;
        RECT 33.330 211.930 33.605 212.100 ;
        RECT 33.325 211.760 33.605 211.930 ;
        RECT 32.610 211.700 32.785 211.735 ;
        RECT 31.855 211.530 32.785 211.700 ;
        RECT 29.585 210.980 30.335 211.500 ;
        RECT 24.820 209.890 25.690 210.230 ;
        RECT 26.280 210.270 27.080 210.440 ;
        RECT 25.860 209.720 26.110 210.180 ;
        RECT 26.280 209.980 26.450 210.270 ;
        RECT 26.630 209.720 26.960 210.100 ;
        RECT 27.255 209.720 27.425 210.780 ;
        RECT 27.635 210.730 29.360 210.900 ;
        RECT 30.505 210.810 31.255 211.330 ;
        RECT 27.635 209.890 27.925 210.730 ;
        RECT 28.095 209.720 28.265 210.560 ;
        RECT 28.475 209.890 28.725 210.730 ;
        RECT 28.935 209.720 29.105 210.560 ;
        RECT 29.585 209.720 31.255 210.810 ;
        RECT 31.430 210.860 31.600 211.530 ;
        RECT 31.855 211.360 32.025 211.530 ;
        RECT 31.770 211.030 32.025 211.360 ;
        RECT 32.250 211.030 32.445 211.360 ;
        RECT 31.430 209.890 31.765 210.860 ;
        RECT 31.935 209.720 32.105 210.860 ;
        RECT 32.275 210.060 32.445 211.030 ;
        RECT 32.615 210.400 32.785 211.530 ;
        RECT 32.955 210.740 33.125 211.540 ;
        RECT 33.330 210.940 33.605 211.760 ;
        RECT 33.775 210.740 33.965 212.100 ;
        RECT 34.145 211.735 34.655 212.270 ;
        RECT 34.875 211.460 35.120 212.065 ;
        RECT 35.575 211.545 35.905 212.055 ;
        RECT 36.075 211.870 36.405 212.270 ;
        RECT 37.455 211.700 37.785 212.040 ;
        RECT 37.955 211.870 38.285 212.270 ;
        RECT 34.165 211.290 35.395 211.460 ;
        RECT 32.955 210.570 33.965 210.740 ;
        RECT 34.135 210.725 34.885 210.915 ;
        RECT 32.615 210.230 33.740 210.400 ;
        RECT 34.135 210.060 34.305 210.725 ;
        RECT 35.055 210.480 35.395 211.290 ;
        RECT 32.275 209.890 34.305 210.060 ;
        RECT 34.475 209.720 34.645 210.480 ;
        RECT 34.880 210.070 35.395 210.480 ;
        RECT 35.575 210.910 35.765 211.545 ;
        RECT 36.075 211.530 38.440 211.700 ;
        RECT 39.705 211.545 39.995 212.270 ;
        RECT 40.625 211.700 41.060 212.100 ;
        RECT 41.230 211.870 41.615 212.270 ;
        RECT 40.625 211.530 41.615 211.700 ;
        RECT 41.785 211.530 42.210 212.100 ;
        RECT 42.400 211.700 42.655 212.100 ;
        RECT 42.825 211.870 43.210 212.270 ;
        RECT 42.400 211.530 43.210 211.700 ;
        RECT 43.380 211.530 43.625 212.100 ;
        RECT 43.815 211.700 44.070 212.100 ;
        RECT 44.240 211.870 44.625 212.270 ;
        RECT 43.815 211.530 44.625 211.700 ;
        RECT 44.795 211.530 45.055 212.100 ;
        RECT 45.285 211.790 45.565 212.270 ;
        RECT 45.735 211.620 45.995 212.010 ;
        RECT 46.170 211.790 46.425 212.270 ;
        RECT 46.595 211.620 46.890 212.010 ;
        RECT 47.070 211.790 47.345 212.270 ;
        RECT 47.515 211.770 47.815 212.100 ;
        RECT 36.075 211.360 36.245 211.530 ;
        RECT 35.935 211.030 36.245 211.360 ;
        RECT 36.415 211.030 36.720 211.360 ;
        RECT 35.575 210.780 35.795 210.910 ;
        RECT 35.575 209.930 35.905 210.780 ;
        RECT 36.075 209.720 36.325 210.860 ;
        RECT 36.505 210.700 36.720 211.030 ;
        RECT 36.895 210.700 37.180 211.360 ;
        RECT 37.375 210.700 37.640 211.360 ;
        RECT 37.855 210.700 38.100 211.360 ;
        RECT 38.270 210.530 38.440 211.530 ;
        RECT 41.280 211.360 41.615 211.530 ;
        RECT 41.860 211.360 42.210 211.530 ;
        RECT 42.860 211.360 43.210 211.530 ;
        RECT 43.455 211.360 43.625 211.530 ;
        RECT 44.275 211.360 44.625 211.530 ;
        RECT 36.515 210.360 37.805 210.530 ;
        RECT 36.515 209.940 36.765 210.360 ;
        RECT 36.995 209.720 37.325 210.190 ;
        RECT 37.555 209.940 37.805 210.360 ;
        RECT 37.985 210.360 38.440 210.530 ;
        RECT 37.985 209.930 38.315 210.360 ;
        RECT 39.705 209.720 39.995 210.885 ;
        RECT 40.625 210.655 41.110 211.360 ;
        RECT 41.280 211.030 41.690 211.360 ;
        RECT 41.280 210.485 41.615 211.030 ;
        RECT 41.860 210.860 42.690 211.360 ;
        RECT 40.625 210.315 41.615 210.485 ;
        RECT 41.785 210.680 42.690 210.860 ;
        RECT 42.860 211.030 43.285 211.360 ;
        RECT 40.625 209.890 41.060 210.315 ;
        RECT 41.230 209.720 41.615 210.145 ;
        RECT 41.785 209.890 42.210 210.680 ;
        RECT 42.860 210.510 43.210 211.030 ;
        RECT 43.455 210.860 44.105 211.360 ;
        RECT 42.380 210.315 43.210 210.510 ;
        RECT 43.380 210.680 44.105 210.860 ;
        RECT 44.275 211.030 44.700 211.360 ;
        RECT 42.380 209.890 42.655 210.315 ;
        RECT 42.825 209.720 43.210 210.145 ;
        RECT 43.380 209.890 43.625 210.680 ;
        RECT 44.275 210.510 44.625 211.030 ;
        RECT 44.870 210.860 45.055 211.530 ;
        RECT 43.815 210.315 44.625 210.510 ;
        RECT 43.815 209.890 44.070 210.315 ;
        RECT 44.240 209.720 44.625 210.145 ;
        RECT 44.795 209.890 45.055 210.860 ;
        RECT 45.240 211.450 46.890 211.620 ;
        RECT 45.240 210.940 45.645 211.450 ;
        RECT 45.815 211.110 46.955 211.280 ;
        RECT 45.240 210.770 45.995 210.940 ;
        RECT 45.280 209.720 45.565 210.590 ;
        RECT 45.735 210.520 45.995 210.770 ;
        RECT 46.785 210.860 46.955 211.110 ;
        RECT 47.125 211.030 47.475 211.600 ;
        RECT 47.645 210.860 47.815 211.770 ;
        RECT 46.785 210.690 47.815 210.860 ;
        RECT 45.735 210.350 46.855 210.520 ;
        RECT 45.735 209.890 45.995 210.350 ;
        RECT 46.170 209.720 46.425 210.180 ;
        RECT 46.595 209.890 46.855 210.350 ;
        RECT 47.025 209.720 47.335 210.520 ;
        RECT 47.505 209.890 47.815 210.690 ;
        RECT 47.985 211.810 48.545 212.100 ;
        RECT 48.715 211.810 48.965 212.270 ;
        RECT 47.985 210.440 48.235 211.810 ;
        RECT 49.585 211.640 49.915 212.000 ;
        RECT 48.525 211.450 49.915 211.640 ;
        RECT 51.205 211.470 51.900 212.100 ;
        RECT 52.105 211.470 52.415 212.270 ;
        RECT 48.525 211.360 48.695 211.450 ;
        RECT 48.405 211.030 48.695 211.360 ;
        RECT 48.865 211.030 49.205 211.280 ;
        RECT 49.425 211.030 50.100 211.280 ;
        RECT 51.225 211.030 51.560 211.280 ;
        RECT 48.525 210.780 48.695 211.030 ;
        RECT 48.525 210.610 49.465 210.780 ;
        RECT 49.835 210.670 50.100 211.030 ;
        RECT 51.730 210.870 51.900 211.470 ;
        RECT 53.050 211.430 53.310 212.270 ;
        RECT 53.485 211.525 53.740 212.100 ;
        RECT 53.910 211.890 54.240 212.270 ;
        RECT 54.455 211.720 54.625 212.100 ;
        RECT 53.910 211.550 54.625 211.720 ;
        RECT 52.070 211.030 52.405 211.300 ;
        RECT 47.985 209.890 48.445 210.440 ;
        RECT 48.635 209.720 48.965 210.440 ;
        RECT 49.165 210.060 49.465 210.610 ;
        RECT 49.635 209.720 49.915 210.390 ;
        RECT 51.205 209.720 51.465 210.860 ;
        RECT 51.635 209.890 51.965 210.870 ;
        RECT 52.135 209.720 52.415 210.860 ;
        RECT 53.050 209.720 53.310 210.870 ;
        RECT 53.485 210.795 53.655 211.525 ;
        RECT 53.910 211.360 54.080 211.550 ;
        RECT 54.890 211.530 55.145 212.100 ;
        RECT 55.315 211.870 55.645 212.270 ;
        RECT 56.070 211.735 56.600 212.100 ;
        RECT 56.070 211.700 56.245 211.735 ;
        RECT 55.315 211.530 56.245 211.700 ;
        RECT 53.825 211.030 54.080 211.360 ;
        RECT 53.910 210.820 54.080 211.030 ;
        RECT 54.360 211.000 54.715 211.370 ;
        RECT 54.890 210.860 55.060 211.530 ;
        RECT 55.315 211.360 55.485 211.530 ;
        RECT 55.230 211.030 55.485 211.360 ;
        RECT 55.710 211.030 55.905 211.360 ;
        RECT 53.485 209.890 53.740 210.795 ;
        RECT 53.910 210.650 54.625 210.820 ;
        RECT 53.910 209.720 54.240 210.480 ;
        RECT 54.455 209.890 54.625 210.650 ;
        RECT 54.890 209.890 55.225 210.860 ;
        RECT 55.395 209.720 55.565 210.860 ;
        RECT 55.735 210.060 55.905 211.030 ;
        RECT 56.075 210.400 56.245 211.530 ;
        RECT 56.415 210.740 56.585 211.540 ;
        RECT 56.790 211.250 57.065 212.100 ;
        RECT 56.785 211.080 57.065 211.250 ;
        RECT 56.790 210.940 57.065 211.080 ;
        RECT 57.235 210.740 57.425 212.100 ;
        RECT 57.605 211.735 58.115 212.270 ;
        RECT 58.335 211.460 58.580 212.065 ;
        RECT 57.625 211.290 58.855 211.460 ;
        RECT 59.085 211.450 59.295 212.270 ;
        RECT 59.465 211.470 59.795 212.100 ;
        RECT 56.415 210.570 57.425 210.740 ;
        RECT 57.595 210.725 58.345 210.915 ;
        RECT 56.075 210.230 57.200 210.400 ;
        RECT 57.595 210.060 57.765 210.725 ;
        RECT 58.515 210.480 58.855 211.290 ;
        RECT 59.465 210.870 59.715 211.470 ;
        RECT 59.965 211.450 60.195 212.270 ;
        RECT 60.680 211.460 60.925 212.065 ;
        RECT 61.145 211.735 61.655 212.270 ;
        RECT 60.405 211.290 61.635 211.460 ;
        RECT 59.885 211.030 60.215 211.280 ;
        RECT 55.735 209.890 57.765 210.060 ;
        RECT 57.935 209.720 58.105 210.480 ;
        RECT 58.340 210.070 58.855 210.480 ;
        RECT 59.085 209.720 59.295 210.860 ;
        RECT 59.465 209.890 59.795 210.870 ;
        RECT 59.965 209.720 60.195 210.860 ;
        RECT 60.405 210.480 60.745 211.290 ;
        RECT 60.915 210.725 61.665 210.915 ;
        RECT 60.405 210.070 60.920 210.480 ;
        RECT 61.155 209.720 61.325 210.480 ;
        RECT 61.495 210.060 61.665 210.725 ;
        RECT 61.835 210.740 62.025 212.100 ;
        RECT 62.195 211.930 62.470 212.100 ;
        RECT 62.195 211.760 62.475 211.930 ;
        RECT 62.195 210.940 62.470 211.760 ;
        RECT 62.660 211.735 63.190 212.100 ;
        RECT 63.615 211.870 63.945 212.270 ;
        RECT 63.015 211.700 63.190 211.735 ;
        RECT 62.675 210.740 62.845 211.540 ;
        RECT 61.835 210.570 62.845 210.740 ;
        RECT 63.015 211.530 63.945 211.700 ;
        RECT 64.115 211.530 64.370 212.100 ;
        RECT 65.465 211.545 65.755 212.270 ;
        RECT 63.015 210.400 63.185 211.530 ;
        RECT 63.775 211.360 63.945 211.530 ;
        RECT 62.060 210.230 63.185 210.400 ;
        RECT 63.355 211.030 63.550 211.360 ;
        RECT 63.775 211.030 64.030 211.360 ;
        RECT 63.355 210.060 63.525 211.030 ;
        RECT 64.200 210.860 64.370 211.530 ;
        RECT 65.925 211.500 68.515 212.270 ;
        RECT 69.150 211.530 69.405 212.100 ;
        RECT 69.575 211.870 69.905 212.270 ;
        RECT 70.330 211.735 70.860 212.100 ;
        RECT 70.330 211.700 70.505 211.735 ;
        RECT 69.575 211.530 70.505 211.700 ;
        RECT 65.925 210.980 67.135 211.500 ;
        RECT 61.495 209.890 63.525 210.060 ;
        RECT 63.695 209.720 63.865 210.860 ;
        RECT 64.035 209.890 64.370 210.860 ;
        RECT 65.465 209.720 65.755 210.885 ;
        RECT 67.305 210.810 68.515 211.330 ;
        RECT 65.925 209.720 68.515 210.810 ;
        RECT 69.150 210.860 69.320 211.530 ;
        RECT 69.575 211.360 69.745 211.530 ;
        RECT 69.490 211.030 69.745 211.360 ;
        RECT 69.970 211.030 70.165 211.360 ;
        RECT 69.150 209.890 69.485 210.860 ;
        RECT 69.655 209.720 69.825 210.860 ;
        RECT 69.995 210.060 70.165 211.030 ;
        RECT 70.335 210.400 70.505 211.530 ;
        RECT 70.675 210.740 70.845 211.540 ;
        RECT 71.050 211.250 71.325 212.100 ;
        RECT 71.045 211.080 71.325 211.250 ;
        RECT 71.050 210.940 71.325 211.080 ;
        RECT 71.495 210.740 71.685 212.100 ;
        RECT 71.865 211.735 72.375 212.270 ;
        RECT 72.595 211.460 72.840 212.065 ;
        RECT 73.285 211.470 73.980 212.100 ;
        RECT 74.185 211.470 74.495 212.270 ;
        RECT 75.585 211.470 76.280 212.100 ;
        RECT 76.485 211.470 76.795 212.270 ;
        RECT 71.885 211.290 73.115 211.460 ;
        RECT 70.675 210.570 71.685 210.740 ;
        RECT 71.855 210.725 72.605 210.915 ;
        RECT 70.335 210.230 71.460 210.400 ;
        RECT 71.855 210.060 72.025 210.725 ;
        RECT 72.775 210.480 73.115 211.290 ;
        RECT 73.305 211.030 73.640 211.280 ;
        RECT 73.810 210.870 73.980 211.470 ;
        RECT 74.150 211.030 74.485 211.300 ;
        RECT 75.605 211.030 75.940 211.280 ;
        RECT 76.110 210.870 76.280 211.470 ;
        RECT 77.700 211.460 77.945 212.065 ;
        RECT 78.165 211.735 78.675 212.270 ;
        RECT 76.450 211.030 76.785 211.300 ;
        RECT 77.425 211.290 78.655 211.460 ;
        RECT 69.995 209.890 72.025 210.060 ;
        RECT 72.195 209.720 72.365 210.480 ;
        RECT 72.600 210.070 73.115 210.480 ;
        RECT 73.285 209.720 73.545 210.860 ;
        RECT 73.715 209.890 74.045 210.870 ;
        RECT 74.215 209.720 74.495 210.860 ;
        RECT 75.585 209.720 75.845 210.860 ;
        RECT 76.015 209.890 76.345 210.870 ;
        RECT 76.515 209.720 76.795 210.860 ;
        RECT 77.425 210.480 77.765 211.290 ;
        RECT 77.935 210.725 78.685 210.915 ;
        RECT 77.425 210.070 77.940 210.480 ;
        RECT 78.175 209.720 78.345 210.480 ;
        RECT 78.515 210.060 78.685 210.725 ;
        RECT 78.855 210.740 79.045 212.100 ;
        RECT 79.215 211.930 79.490 212.100 ;
        RECT 79.215 211.760 79.495 211.930 ;
        RECT 79.215 210.940 79.490 211.760 ;
        RECT 79.680 211.735 80.210 212.100 ;
        RECT 80.635 211.870 80.965 212.270 ;
        RECT 80.035 211.700 80.210 211.735 ;
        RECT 79.695 210.740 79.865 211.540 ;
        RECT 78.855 210.570 79.865 210.740 ;
        RECT 80.035 211.530 80.965 211.700 ;
        RECT 81.135 211.530 81.390 212.100 ;
        RECT 80.035 210.400 80.205 211.530 ;
        RECT 80.795 211.360 80.965 211.530 ;
        RECT 79.080 210.230 80.205 210.400 ;
        RECT 80.375 211.030 80.570 211.360 ;
        RECT 80.795 211.030 81.050 211.360 ;
        RECT 80.375 210.060 80.545 211.030 ;
        RECT 81.220 210.860 81.390 211.530 ;
        RECT 78.515 209.890 80.545 210.060 ;
        RECT 80.715 209.720 80.885 210.860 ;
        RECT 81.055 209.890 81.390 210.860 ;
        RECT 81.565 211.770 81.825 212.100 ;
        RECT 82.035 211.790 82.310 212.270 ;
        RECT 81.565 210.860 81.735 211.770 ;
        RECT 82.520 211.700 82.725 212.100 ;
        RECT 82.895 211.870 83.230 212.270 ;
        RECT 81.905 211.030 82.265 211.610 ;
        RECT 82.520 211.530 83.205 211.700 ;
        RECT 82.445 210.860 82.695 211.360 ;
        RECT 81.565 210.690 82.695 210.860 ;
        RECT 81.565 209.920 81.835 210.690 ;
        RECT 82.865 210.500 83.205 211.530 ;
        RECT 83.465 211.450 83.675 212.270 ;
        RECT 83.845 211.470 84.175 212.100 ;
        RECT 83.845 210.870 84.095 211.470 ;
        RECT 84.345 211.450 84.575 212.270 ;
        RECT 85.520 211.460 85.765 212.065 ;
        RECT 85.985 211.735 86.495 212.270 ;
        RECT 85.245 211.290 86.475 211.460 ;
        RECT 84.265 211.030 84.595 211.280 ;
        RECT 82.005 209.720 82.335 210.500 ;
        RECT 82.540 210.325 83.205 210.500 ;
        RECT 82.540 209.920 82.725 210.325 ;
        RECT 82.895 209.720 83.230 210.145 ;
        RECT 83.465 209.720 83.675 210.860 ;
        RECT 83.845 209.890 84.175 210.870 ;
        RECT 84.345 209.720 84.575 210.860 ;
        RECT 85.245 210.480 85.585 211.290 ;
        RECT 85.755 210.725 86.505 210.915 ;
        RECT 85.245 210.070 85.760 210.480 ;
        RECT 85.995 209.720 86.165 210.480 ;
        RECT 86.335 210.060 86.505 210.725 ;
        RECT 86.675 210.740 86.865 212.100 ;
        RECT 87.035 211.930 87.310 212.100 ;
        RECT 87.035 211.760 87.315 211.930 ;
        RECT 87.035 210.940 87.310 211.760 ;
        RECT 87.500 211.735 88.030 212.100 ;
        RECT 88.455 211.870 88.785 212.270 ;
        RECT 87.855 211.700 88.030 211.735 ;
        RECT 87.515 210.740 87.685 211.540 ;
        RECT 86.675 210.570 87.685 210.740 ;
        RECT 87.855 211.530 88.785 211.700 ;
        RECT 88.955 211.530 89.210 212.100 ;
        RECT 87.855 210.400 88.025 211.530 ;
        RECT 88.615 211.360 88.785 211.530 ;
        RECT 86.900 210.230 88.025 210.400 ;
        RECT 88.195 211.030 88.390 211.360 ;
        RECT 88.615 211.030 88.870 211.360 ;
        RECT 88.195 210.060 88.365 211.030 ;
        RECT 89.040 210.860 89.210 211.530 ;
        RECT 89.385 211.470 89.695 212.270 ;
        RECT 89.900 211.470 90.595 212.100 ;
        RECT 91.225 211.545 91.515 212.270 ;
        RECT 91.695 211.910 93.765 212.100 ;
        RECT 93.995 211.910 94.325 212.270 ;
        RECT 94.855 211.910 95.185 212.270 ;
        RECT 95.715 211.910 96.045 212.270 ;
        RECT 92.645 211.890 93.765 211.910 ;
        RECT 89.395 211.030 89.730 211.300 ;
        RECT 89.900 210.870 90.070 211.470 ;
        RECT 90.240 211.030 90.575 211.280 ;
        RECT 86.335 209.890 88.365 210.060 ;
        RECT 88.535 209.720 88.705 210.860 ;
        RECT 88.875 209.890 89.210 210.860 ;
        RECT 89.385 209.720 89.665 210.860 ;
        RECT 89.835 209.890 90.165 210.870 ;
        RECT 90.335 209.720 90.595 210.860 ;
        RECT 91.225 209.720 91.515 210.885 ;
        RECT 91.685 210.385 91.975 211.360 ;
        RECT 92.145 210.815 92.475 211.685 ;
        RECT 92.645 211.465 92.835 211.890 ;
        RECT 96.290 211.870 96.625 212.270 ;
        RECT 95.355 211.720 95.545 211.840 ;
        RECT 93.005 211.510 95.545 211.720 ;
        RECT 96.795 211.700 97.000 212.100 ;
        RECT 97.210 211.790 97.485 212.270 ;
        RECT 97.695 211.770 97.955 212.100 ;
        RECT 95.715 211.280 96.055 211.590 ;
        RECT 92.645 210.990 93.505 211.280 ;
        RECT 93.965 211.000 94.935 211.280 ;
        RECT 95.105 211.110 96.055 211.280 ;
        RECT 95.160 211.060 96.055 211.110 ;
        RECT 96.315 211.530 97.000 211.700 ;
        RECT 92.145 210.645 94.755 210.815 ;
        RECT 91.715 209.720 91.975 210.180 ;
        RECT 92.145 209.890 92.405 210.645 ;
        RECT 92.575 209.720 92.905 210.440 ;
        RECT 93.075 209.890 93.265 210.645 ;
        RECT 93.435 209.720 93.765 210.440 ;
        RECT 93.995 210.060 94.255 210.255 ;
        RECT 94.425 210.230 94.755 210.645 ;
        RECT 94.925 210.660 96.045 210.830 ;
        RECT 94.925 210.060 95.115 210.660 ;
        RECT 93.995 209.890 95.115 210.060 ;
        RECT 95.285 209.720 95.615 210.490 ;
        RECT 95.785 209.890 96.045 210.660 ;
        RECT 96.315 210.500 96.655 211.530 ;
        RECT 96.825 210.860 97.075 211.360 ;
        RECT 97.255 211.030 97.615 211.610 ;
        RECT 97.785 210.860 97.955 211.770 ;
        RECT 98.590 211.720 98.845 212.010 ;
        RECT 99.015 211.890 99.345 212.270 ;
        RECT 98.590 211.550 99.340 211.720 ;
        RECT 96.825 210.690 97.955 210.860 ;
        RECT 98.590 210.730 98.940 211.380 ;
        RECT 96.315 210.325 96.980 210.500 ;
        RECT 96.290 209.720 96.625 210.145 ;
        RECT 96.795 209.920 96.980 210.325 ;
        RECT 97.185 209.720 97.515 210.500 ;
        RECT 97.685 209.920 97.955 210.690 ;
        RECT 99.110 210.560 99.340 211.550 ;
        RECT 98.590 210.390 99.340 210.560 ;
        RECT 98.590 209.890 98.845 210.390 ;
        RECT 99.015 209.720 99.345 210.220 ;
        RECT 99.515 209.890 99.685 212.010 ;
        RECT 100.045 211.910 100.375 212.270 ;
        RECT 100.545 211.880 101.040 212.050 ;
        RECT 101.245 211.880 102.100 212.050 ;
        RECT 99.915 210.690 100.375 211.740 ;
        RECT 99.855 209.905 100.180 210.690 ;
        RECT 100.545 210.520 100.715 211.880 ;
        RECT 100.885 210.970 101.235 211.590 ;
        RECT 101.405 211.370 101.760 211.590 ;
        RECT 101.405 210.780 101.575 211.370 ;
        RECT 101.930 211.170 102.100 211.880 ;
        RECT 102.975 211.810 103.305 212.270 ;
        RECT 103.515 211.910 103.865 212.080 ;
        RECT 102.305 211.340 103.095 211.590 ;
        RECT 103.515 211.520 103.775 211.910 ;
        RECT 104.085 211.820 105.035 212.100 ;
        RECT 105.205 211.830 105.395 212.270 ;
        RECT 105.565 211.890 106.635 212.060 ;
        RECT 103.265 211.170 103.435 211.350 ;
        RECT 100.545 210.350 100.940 210.520 ;
        RECT 101.110 210.390 101.575 210.780 ;
        RECT 101.745 211.000 103.435 211.170 ;
        RECT 100.770 210.220 100.940 210.350 ;
        RECT 101.745 210.220 101.915 211.000 ;
        RECT 103.605 210.830 103.775 211.520 ;
        RECT 102.275 210.660 103.775 210.830 ;
        RECT 103.965 210.860 104.175 211.650 ;
        RECT 104.345 211.030 104.695 211.650 ;
        RECT 104.865 211.040 105.035 211.820 ;
        RECT 105.565 211.660 105.735 211.890 ;
        RECT 105.205 211.490 105.735 211.660 ;
        RECT 105.205 211.210 105.425 211.490 ;
        RECT 105.905 211.320 106.145 211.720 ;
        RECT 104.865 210.870 105.270 211.040 ;
        RECT 105.605 210.950 106.145 211.320 ;
        RECT 106.315 211.535 106.635 211.890 ;
        RECT 106.880 211.810 107.185 212.270 ;
        RECT 107.355 211.560 107.610 212.090 ;
        RECT 107.785 211.760 108.090 212.270 ;
        RECT 106.315 211.360 106.640 211.535 ;
        RECT 106.315 211.060 107.230 211.360 ;
        RECT 106.490 211.030 107.230 211.060 ;
        RECT 103.965 210.700 104.640 210.860 ;
        RECT 105.100 210.780 105.270 210.870 ;
        RECT 103.965 210.690 104.930 210.700 ;
        RECT 103.605 210.520 103.775 210.660 ;
        RECT 100.350 209.720 100.600 210.180 ;
        RECT 100.770 209.890 101.020 210.220 ;
        RECT 101.235 209.890 101.915 210.220 ;
        RECT 102.085 210.320 103.160 210.490 ;
        RECT 103.605 210.350 104.165 210.520 ;
        RECT 104.470 210.400 104.930 210.690 ;
        RECT 105.100 210.610 106.320 210.780 ;
        RECT 102.085 209.980 102.255 210.320 ;
        RECT 102.490 209.720 102.820 210.150 ;
        RECT 102.990 209.980 103.160 210.320 ;
        RECT 103.455 209.720 103.825 210.180 ;
        RECT 103.995 209.890 104.165 210.350 ;
        RECT 105.100 210.230 105.270 210.610 ;
        RECT 106.490 210.440 106.660 211.030 ;
        RECT 107.400 210.910 107.610 211.560 ;
        RECT 107.785 211.030 108.100 211.590 ;
        RECT 108.270 211.280 108.520 212.090 ;
        RECT 108.690 211.745 108.950 212.270 ;
        RECT 109.130 211.280 109.380 212.090 ;
        RECT 109.550 211.710 109.810 212.270 ;
        RECT 109.980 211.620 110.240 212.075 ;
        RECT 110.410 211.790 110.670 212.270 ;
        RECT 110.840 211.620 111.100 212.075 ;
        RECT 111.270 211.790 111.530 212.270 ;
        RECT 111.700 211.620 111.960 212.075 ;
        RECT 112.130 211.790 112.375 212.270 ;
        RECT 112.545 211.620 112.820 212.075 ;
        RECT 112.990 211.790 113.235 212.270 ;
        RECT 113.405 211.620 113.665 212.075 ;
        RECT 113.845 211.790 114.095 212.270 ;
        RECT 114.265 211.620 114.525 212.075 ;
        RECT 114.705 211.790 114.955 212.270 ;
        RECT 115.125 211.620 115.385 212.075 ;
        RECT 115.565 211.790 115.825 212.270 ;
        RECT 115.995 211.620 116.255 212.075 ;
        RECT 116.425 211.790 116.725 212.270 ;
        RECT 109.980 211.450 116.725 211.620 ;
        RECT 116.985 211.545 117.275 212.270 ;
        RECT 117.450 211.870 117.785 212.270 ;
        RECT 117.955 211.700 118.160 212.100 ;
        RECT 118.370 211.790 118.645 212.270 ;
        RECT 118.855 211.770 119.115 212.100 ;
        RECT 119.615 211.870 119.945 212.270 ;
        RECT 108.270 211.030 115.390 211.280 ;
        RECT 104.400 209.890 105.270 210.230 ;
        RECT 105.860 210.270 106.660 210.440 ;
        RECT 105.440 209.720 105.690 210.180 ;
        RECT 105.860 209.980 106.030 210.270 ;
        RECT 106.210 209.720 106.540 210.100 ;
        RECT 106.880 209.720 107.185 210.860 ;
        RECT 107.355 210.030 107.610 210.910 ;
        RECT 107.795 209.720 108.090 210.530 ;
        RECT 108.270 209.890 108.515 211.030 ;
        RECT 108.690 209.720 108.950 210.530 ;
        RECT 109.130 209.895 109.380 211.030 ;
        RECT 115.560 210.910 116.725 211.450 ;
        RECT 117.475 211.530 118.160 211.700 ;
        RECT 115.560 210.860 116.755 210.910 ;
        RECT 109.980 210.740 116.755 210.860 ;
        RECT 109.980 210.635 116.725 210.740 ;
        RECT 109.980 210.620 115.385 210.635 ;
        RECT 109.550 209.725 109.810 210.520 ;
        RECT 109.980 209.895 110.240 210.620 ;
        RECT 110.410 209.725 110.670 210.450 ;
        RECT 110.840 209.895 111.100 210.620 ;
        RECT 111.270 209.725 111.530 210.450 ;
        RECT 111.700 209.895 111.960 210.620 ;
        RECT 112.130 209.725 112.390 210.450 ;
        RECT 112.560 209.895 112.820 210.620 ;
        RECT 112.990 209.725 113.235 210.450 ;
        RECT 113.405 209.895 113.665 210.620 ;
        RECT 113.850 209.725 114.095 210.450 ;
        RECT 114.265 209.895 114.525 210.620 ;
        RECT 114.710 209.725 114.955 210.450 ;
        RECT 115.125 209.895 115.385 210.620 ;
        RECT 115.570 209.725 115.825 210.450 ;
        RECT 115.995 209.895 116.285 210.635 ;
        RECT 109.550 209.720 115.825 209.725 ;
        RECT 116.455 209.720 116.725 210.465 ;
        RECT 116.985 209.720 117.275 210.885 ;
        RECT 117.475 210.500 117.815 211.530 ;
        RECT 117.985 210.860 118.235 211.360 ;
        RECT 118.415 211.030 118.775 211.610 ;
        RECT 118.945 210.860 119.115 211.770 ;
        RECT 120.115 211.700 120.445 212.040 ;
        RECT 121.495 211.870 121.825 212.270 ;
        RECT 117.985 210.690 119.115 210.860 ;
        RECT 117.475 210.325 118.140 210.500 ;
        RECT 117.450 209.720 117.785 210.145 ;
        RECT 117.955 209.920 118.140 210.325 ;
        RECT 118.345 209.720 118.675 210.500 ;
        RECT 118.845 209.920 119.115 210.690 ;
        RECT 119.460 211.530 121.825 211.700 ;
        RECT 121.995 211.545 122.325 212.055 ;
        RECT 119.460 210.530 119.630 211.530 ;
        RECT 121.655 211.360 121.825 211.530 ;
        RECT 119.800 210.700 120.045 211.360 ;
        RECT 120.260 210.700 120.525 211.360 ;
        RECT 120.720 210.700 121.005 211.360 ;
        RECT 121.180 211.030 121.485 211.360 ;
        RECT 121.655 211.030 121.965 211.360 ;
        RECT 121.180 210.700 121.395 211.030 ;
        RECT 119.460 210.360 119.915 210.530 ;
        RECT 119.585 209.930 119.915 210.360 ;
        RECT 120.095 210.360 121.385 210.530 ;
        RECT 120.095 209.940 120.345 210.360 ;
        RECT 120.575 209.720 120.905 210.190 ;
        RECT 121.135 209.940 121.385 210.360 ;
        RECT 121.575 209.720 121.825 210.860 ;
        RECT 122.135 210.780 122.325 211.545 ;
        RECT 122.565 211.450 122.775 212.270 ;
        RECT 122.945 211.470 123.275 212.100 ;
        RECT 122.945 210.870 123.195 211.470 ;
        RECT 123.445 211.450 123.675 212.270 ;
        RECT 123.890 211.720 124.145 212.010 ;
        RECT 124.315 211.890 124.645 212.270 ;
        RECT 123.890 211.550 124.640 211.720 ;
        RECT 123.365 211.030 123.695 211.280 ;
        RECT 121.995 209.930 122.325 210.780 ;
        RECT 122.565 209.720 122.775 210.860 ;
        RECT 122.945 209.890 123.275 210.870 ;
        RECT 123.445 209.720 123.675 210.860 ;
        RECT 123.890 210.730 124.240 211.380 ;
        RECT 124.410 210.560 124.640 211.550 ;
        RECT 123.890 210.390 124.640 210.560 ;
        RECT 123.890 209.890 124.145 210.390 ;
        RECT 124.315 209.720 124.645 210.220 ;
        RECT 124.815 209.890 124.985 212.010 ;
        RECT 125.345 211.910 125.675 212.270 ;
        RECT 125.845 211.880 126.340 212.050 ;
        RECT 126.545 211.880 127.400 212.050 ;
        RECT 125.215 210.690 125.675 211.740 ;
        RECT 125.155 209.905 125.480 210.690 ;
        RECT 125.845 210.520 126.015 211.880 ;
        RECT 126.185 210.970 126.535 211.590 ;
        RECT 126.705 211.370 127.060 211.590 ;
        RECT 126.705 210.780 126.875 211.370 ;
        RECT 127.230 211.170 127.400 211.880 ;
        RECT 128.275 211.810 128.605 212.270 ;
        RECT 128.815 211.910 129.165 212.080 ;
        RECT 127.605 211.340 128.395 211.590 ;
        RECT 128.815 211.520 129.075 211.910 ;
        RECT 129.385 211.820 130.335 212.100 ;
        RECT 130.505 211.830 130.695 212.270 ;
        RECT 130.865 211.890 131.935 212.060 ;
        RECT 128.565 211.170 128.735 211.350 ;
        RECT 125.845 210.350 126.240 210.520 ;
        RECT 126.410 210.390 126.875 210.780 ;
        RECT 127.045 211.000 128.735 211.170 ;
        RECT 126.070 210.220 126.240 210.350 ;
        RECT 127.045 210.220 127.215 211.000 ;
        RECT 128.905 210.830 129.075 211.520 ;
        RECT 127.575 210.660 129.075 210.830 ;
        RECT 129.265 210.860 129.475 211.650 ;
        RECT 129.645 211.030 129.995 211.650 ;
        RECT 130.165 211.040 130.335 211.820 ;
        RECT 130.865 211.660 131.035 211.890 ;
        RECT 130.505 211.490 131.035 211.660 ;
        RECT 130.505 211.210 130.725 211.490 ;
        RECT 131.205 211.320 131.445 211.720 ;
        RECT 130.165 210.870 130.570 211.040 ;
        RECT 130.905 210.950 131.445 211.320 ;
        RECT 131.615 211.535 131.935 211.890 ;
        RECT 132.180 211.810 132.485 212.270 ;
        RECT 132.655 211.560 132.910 212.090 ;
        RECT 131.615 211.360 131.940 211.535 ;
        RECT 131.615 211.060 132.530 211.360 ;
        RECT 131.790 211.030 132.530 211.060 ;
        RECT 129.265 210.700 129.940 210.860 ;
        RECT 130.400 210.780 130.570 210.870 ;
        RECT 129.265 210.690 130.230 210.700 ;
        RECT 128.905 210.520 129.075 210.660 ;
        RECT 125.650 209.720 125.900 210.180 ;
        RECT 126.070 209.890 126.320 210.220 ;
        RECT 126.535 209.890 127.215 210.220 ;
        RECT 127.385 210.320 128.460 210.490 ;
        RECT 128.905 210.350 129.465 210.520 ;
        RECT 129.770 210.400 130.230 210.690 ;
        RECT 130.400 210.610 131.620 210.780 ;
        RECT 127.385 209.980 127.555 210.320 ;
        RECT 127.790 209.720 128.120 210.150 ;
        RECT 128.290 209.980 128.460 210.320 ;
        RECT 128.755 209.720 129.125 210.180 ;
        RECT 129.295 209.890 129.465 210.350 ;
        RECT 130.400 210.230 130.570 210.610 ;
        RECT 131.790 210.440 131.960 211.030 ;
        RECT 132.700 210.910 132.910 211.560 ;
        RECT 129.700 209.890 130.570 210.230 ;
        RECT 131.160 210.270 131.960 210.440 ;
        RECT 130.740 209.720 130.990 210.180 ;
        RECT 131.160 209.980 131.330 210.270 ;
        RECT 131.510 209.720 131.840 210.100 ;
        RECT 132.180 209.720 132.485 210.860 ;
        RECT 132.655 210.030 132.910 210.910 ;
        RECT 133.090 211.530 133.345 212.100 ;
        RECT 133.515 211.870 133.845 212.270 ;
        RECT 134.270 211.735 134.800 212.100 ;
        RECT 134.270 211.700 134.445 211.735 ;
        RECT 133.515 211.530 134.445 211.700 ;
        RECT 134.990 211.590 135.265 212.100 ;
        RECT 133.090 210.860 133.260 211.530 ;
        RECT 133.515 211.360 133.685 211.530 ;
        RECT 133.430 211.030 133.685 211.360 ;
        RECT 133.910 211.030 134.105 211.360 ;
        RECT 133.090 209.890 133.425 210.860 ;
        RECT 133.595 209.720 133.765 210.860 ;
        RECT 133.935 210.060 134.105 211.030 ;
        RECT 134.275 210.400 134.445 211.530 ;
        RECT 134.615 210.740 134.785 211.540 ;
        RECT 134.985 211.420 135.265 211.590 ;
        RECT 134.990 210.940 135.265 211.420 ;
        RECT 135.435 210.740 135.625 212.100 ;
        RECT 135.805 211.735 136.315 212.270 ;
        RECT 136.535 211.460 136.780 212.065 ;
        RECT 137.225 211.500 140.735 212.270 ;
        RECT 140.995 211.720 141.165 212.100 ;
        RECT 141.380 211.890 141.710 212.270 ;
        RECT 140.995 211.550 141.710 211.720 ;
        RECT 135.825 211.290 137.055 211.460 ;
        RECT 134.615 210.570 135.625 210.740 ;
        RECT 135.795 210.725 136.545 210.915 ;
        RECT 134.275 210.230 135.400 210.400 ;
        RECT 135.795 210.060 135.965 210.725 ;
        RECT 136.715 210.480 137.055 211.290 ;
        RECT 137.225 210.980 138.875 211.500 ;
        RECT 139.045 210.810 140.735 211.330 ;
        RECT 140.905 211.000 141.260 211.370 ;
        RECT 141.540 211.360 141.710 211.550 ;
        RECT 141.880 211.525 142.135 212.100 ;
        RECT 141.540 211.030 141.795 211.360 ;
        RECT 141.540 210.820 141.710 211.030 ;
        RECT 133.935 209.890 135.965 210.060 ;
        RECT 136.135 209.720 136.305 210.480 ;
        RECT 136.540 210.070 137.055 210.480 ;
        RECT 137.225 209.720 140.735 210.810 ;
        RECT 140.995 210.650 141.710 210.820 ;
        RECT 141.965 210.795 142.135 211.525 ;
        RECT 142.310 211.430 142.570 212.270 ;
        RECT 142.745 211.545 143.035 212.270 ;
        RECT 143.205 211.520 144.415 212.270 ;
        RECT 144.675 211.720 144.845 212.100 ;
        RECT 145.060 211.890 145.390 212.270 ;
        RECT 144.675 211.550 145.390 211.720 ;
        RECT 143.205 210.980 143.725 211.520 ;
        RECT 140.995 209.890 141.165 210.650 ;
        RECT 141.380 209.720 141.710 210.480 ;
        RECT 141.880 209.890 142.135 210.795 ;
        RECT 142.310 209.720 142.570 210.870 ;
        RECT 142.745 209.720 143.035 210.885 ;
        RECT 143.895 210.810 144.415 211.350 ;
        RECT 144.585 211.000 144.940 211.370 ;
        RECT 145.220 211.360 145.390 211.550 ;
        RECT 145.560 211.525 145.815 212.100 ;
        RECT 145.220 211.030 145.475 211.360 ;
        RECT 145.220 210.820 145.390 211.030 ;
        RECT 143.205 209.720 144.415 210.810 ;
        RECT 144.675 210.650 145.390 210.820 ;
        RECT 145.645 210.795 145.815 211.525 ;
        RECT 145.990 211.430 146.250 212.270 ;
        RECT 146.425 211.520 147.635 212.270 ;
        RECT 144.675 209.890 144.845 210.650 ;
        RECT 145.060 209.720 145.390 210.480 ;
        RECT 145.560 209.890 145.815 210.795 ;
        RECT 145.990 209.720 146.250 210.870 ;
        RECT 146.425 210.810 146.945 211.350 ;
        RECT 147.115 210.980 147.635 211.520 ;
        RECT 146.425 209.720 147.635 210.810 ;
        RECT 13.860 209.550 147.720 209.720 ;
        RECT 13.945 208.460 15.155 209.550 ;
        RECT 13.945 207.750 14.465 208.290 ;
        RECT 14.635 207.920 15.155 208.460 ;
        RECT 15.330 208.400 15.590 209.550 ;
        RECT 15.765 208.475 16.020 209.380 ;
        RECT 16.190 208.790 16.520 209.550 ;
        RECT 16.735 208.620 16.905 209.380 ;
        RECT 13.945 207.000 15.155 207.750 ;
        RECT 15.330 207.000 15.590 207.840 ;
        RECT 15.765 207.745 15.935 208.475 ;
        RECT 16.190 208.450 16.905 208.620 ;
        RECT 16.190 208.240 16.360 208.450 ;
        RECT 17.170 208.400 17.430 209.550 ;
        RECT 17.605 208.475 17.860 209.380 ;
        RECT 18.030 208.790 18.360 209.550 ;
        RECT 18.575 208.620 18.745 209.380 ;
        RECT 16.105 207.910 16.360 208.240 ;
        RECT 15.765 207.170 16.020 207.745 ;
        RECT 16.190 207.720 16.360 207.910 ;
        RECT 16.640 207.900 16.995 208.270 ;
        RECT 16.190 207.550 16.905 207.720 ;
        RECT 16.190 207.000 16.520 207.380 ;
        RECT 16.735 207.170 16.905 207.550 ;
        RECT 17.170 207.000 17.430 207.840 ;
        RECT 17.605 207.745 17.775 208.475 ;
        RECT 18.030 208.450 18.745 208.620 ;
        RECT 19.005 208.460 22.515 209.550 ;
        RECT 22.685 208.460 23.895 209.550 ;
        RECT 18.030 208.240 18.200 208.450 ;
        RECT 17.945 207.910 18.200 208.240 ;
        RECT 17.605 207.170 17.860 207.745 ;
        RECT 18.030 207.720 18.200 207.910 ;
        RECT 18.480 207.900 18.835 208.270 ;
        RECT 19.005 207.770 20.655 208.290 ;
        RECT 20.825 207.940 22.515 208.460 ;
        RECT 18.030 207.550 18.745 207.720 ;
        RECT 18.030 207.000 18.360 207.380 ;
        RECT 18.575 207.170 18.745 207.550 ;
        RECT 19.005 207.000 22.515 207.770 ;
        RECT 22.685 207.750 23.205 208.290 ;
        RECT 23.375 207.920 23.895 208.460 ;
        RECT 24.065 208.580 24.655 209.380 ;
        RECT 24.825 208.750 25.110 209.550 ;
        RECT 25.280 208.580 25.610 209.380 ;
        RECT 24.065 208.410 25.610 208.580 ;
        RECT 25.780 208.410 26.030 209.550 ;
        RECT 26.230 208.510 26.655 208.840 ;
        RECT 22.685 207.000 23.895 207.750 ;
        RECT 24.065 207.400 24.355 208.410 ;
        RECT 24.525 207.740 24.695 208.240 ;
        RECT 24.985 207.910 25.315 208.240 ;
        RECT 25.505 207.910 25.775 208.240 ;
        RECT 25.965 207.910 26.315 208.240 ;
        RECT 26.485 207.740 26.655 208.510 ;
        RECT 26.825 208.385 27.115 209.550 ;
        RECT 27.290 208.410 27.625 209.380 ;
        RECT 27.795 208.410 27.965 209.550 ;
        RECT 28.135 209.210 30.165 209.380 ;
        RECT 24.525 207.570 26.655 207.740 ;
        RECT 27.290 207.740 27.460 208.410 ;
        RECT 28.135 208.240 28.305 209.210 ;
        RECT 27.630 207.910 27.885 208.240 ;
        RECT 28.110 207.910 28.305 208.240 ;
        RECT 28.475 208.870 29.600 209.040 ;
        RECT 27.715 207.740 27.885 207.910 ;
        RECT 28.475 207.740 28.645 208.870 ;
        RECT 24.065 207.170 24.655 207.400 ;
        RECT 25.700 207.000 26.030 207.400 ;
        RECT 26.230 207.360 26.655 207.570 ;
        RECT 26.825 207.000 27.115 207.725 ;
        RECT 27.290 207.170 27.545 207.740 ;
        RECT 27.715 207.570 28.645 207.740 ;
        RECT 28.815 208.530 29.825 208.700 ;
        RECT 28.815 207.730 28.985 208.530 ;
        RECT 29.190 208.190 29.465 208.330 ;
        RECT 29.185 208.020 29.465 208.190 ;
        RECT 28.470 207.535 28.645 207.570 ;
        RECT 27.715 207.000 28.045 207.400 ;
        RECT 28.470 207.170 29.000 207.535 ;
        RECT 29.190 207.170 29.465 208.020 ;
        RECT 29.635 207.170 29.825 208.530 ;
        RECT 29.995 208.545 30.165 209.210 ;
        RECT 30.335 208.790 30.505 209.550 ;
        RECT 30.740 208.790 31.255 209.200 ;
        RECT 29.995 208.355 30.745 208.545 ;
        RECT 30.915 207.980 31.255 208.790 ;
        RECT 30.025 207.810 31.255 207.980 ;
        RECT 31.435 208.490 31.765 209.340 ;
        RECT 31.435 208.360 31.655 208.490 ;
        RECT 31.935 208.410 32.185 209.550 ;
        RECT 32.375 208.910 32.625 209.330 ;
        RECT 32.855 209.080 33.185 209.550 ;
        RECT 33.415 208.910 33.665 209.330 ;
        RECT 32.375 208.740 33.665 208.910 ;
        RECT 33.845 208.910 34.175 209.340 ;
        RECT 33.845 208.740 34.300 208.910 ;
        RECT 30.005 207.000 30.515 207.535 ;
        RECT 30.735 207.205 30.980 207.810 ;
        RECT 31.435 207.725 31.625 208.360 ;
        RECT 32.365 208.240 32.580 208.570 ;
        RECT 31.795 207.910 32.105 208.240 ;
        RECT 32.275 207.910 32.580 208.240 ;
        RECT 32.755 207.910 33.040 208.570 ;
        RECT 33.235 207.910 33.500 208.570 ;
        RECT 33.715 207.910 33.960 208.570 ;
        RECT 31.935 207.740 32.105 207.910 ;
        RECT 34.130 207.740 34.300 208.740 ;
        RECT 31.435 207.215 31.765 207.725 ;
        RECT 31.935 207.570 34.300 207.740 ;
        RECT 34.645 208.510 35.070 208.840 ;
        RECT 34.645 207.740 34.815 208.510 ;
        RECT 35.270 208.410 35.520 209.550 ;
        RECT 35.690 208.580 36.020 209.380 ;
        RECT 36.190 208.750 36.475 209.550 ;
        RECT 36.645 208.580 37.235 209.380 ;
        RECT 35.690 208.410 37.235 208.580 ;
        RECT 37.405 208.410 37.685 209.550 ;
        RECT 34.985 207.910 35.335 208.240 ;
        RECT 35.525 207.910 35.795 208.240 ;
        RECT 35.985 207.910 36.315 208.240 ;
        RECT 36.605 207.740 36.775 208.240 ;
        RECT 34.645 207.570 36.775 207.740 ;
        RECT 31.935 207.000 32.265 207.400 ;
        RECT 33.315 207.230 33.645 207.570 ;
        RECT 33.815 207.000 34.145 207.400 ;
        RECT 34.645 207.360 35.070 207.570 ;
        RECT 36.945 207.400 37.235 208.410 ;
        RECT 37.855 208.400 38.185 209.380 ;
        RECT 38.355 208.410 38.615 209.550 ;
        RECT 38.790 208.410 39.125 209.380 ;
        RECT 39.295 208.410 39.465 209.550 ;
        RECT 39.635 209.210 41.665 209.380 ;
        RECT 37.415 207.970 37.750 208.240 ;
        RECT 37.920 207.800 38.090 208.400 ;
        RECT 38.260 207.990 38.595 208.240 ;
        RECT 35.270 207.000 35.600 207.400 ;
        RECT 36.645 207.170 37.235 207.400 ;
        RECT 37.405 207.000 37.715 207.800 ;
        RECT 37.920 207.170 38.615 207.800 ;
        RECT 38.790 207.740 38.960 208.410 ;
        RECT 39.635 208.240 39.805 209.210 ;
        RECT 39.130 207.910 39.385 208.240 ;
        RECT 39.610 207.910 39.805 208.240 ;
        RECT 39.975 208.870 41.100 209.040 ;
        RECT 39.215 207.740 39.385 207.910 ;
        RECT 39.975 207.740 40.145 208.870 ;
        RECT 38.790 207.170 39.045 207.740 ;
        RECT 39.215 207.570 40.145 207.740 ;
        RECT 40.315 208.530 41.325 208.700 ;
        RECT 40.315 207.730 40.485 208.530 ;
        RECT 39.970 207.535 40.145 207.570 ;
        RECT 39.215 207.000 39.545 207.400 ;
        RECT 39.970 207.170 40.500 207.535 ;
        RECT 40.690 207.510 40.965 208.330 ;
        RECT 40.685 207.340 40.965 207.510 ;
        RECT 40.690 207.170 40.965 207.340 ;
        RECT 41.135 207.170 41.325 208.530 ;
        RECT 41.495 208.545 41.665 209.210 ;
        RECT 41.835 208.790 42.005 209.550 ;
        RECT 42.240 208.790 42.755 209.200 ;
        RECT 41.495 208.355 42.245 208.545 ;
        RECT 42.415 207.980 42.755 208.790 ;
        RECT 42.965 208.410 43.195 209.550 ;
        RECT 43.365 208.400 43.695 209.380 ;
        RECT 43.865 208.410 44.075 209.550 ;
        RECT 42.945 207.990 43.275 208.240 ;
        RECT 41.525 207.810 42.755 207.980 ;
        RECT 41.505 207.000 42.015 207.535 ;
        RECT 42.235 207.205 42.480 207.810 ;
        RECT 42.965 207.000 43.195 207.820 ;
        RECT 43.445 207.800 43.695 208.400 ;
        RECT 43.365 207.170 43.695 207.800 ;
        RECT 43.865 207.000 44.075 207.820 ;
        RECT 44.315 207.180 44.575 209.370 ;
        RECT 44.745 208.820 45.085 209.550 ;
        RECT 45.265 208.640 45.535 209.370 ;
        RECT 44.765 208.420 45.535 208.640 ;
        RECT 45.715 208.660 45.945 209.370 ;
        RECT 46.115 208.840 46.445 209.550 ;
        RECT 46.615 208.660 46.875 209.370 ;
        RECT 45.715 208.420 46.875 208.660 ;
        RECT 44.765 207.750 45.055 208.420 ;
        RECT 47.065 208.410 47.340 209.380 ;
        RECT 47.550 208.750 47.830 209.550 ;
        RECT 48.000 209.040 49.615 209.370 ;
        RECT 48.000 208.700 49.175 208.870 ;
        RECT 48.000 208.580 48.170 208.700 ;
        RECT 47.510 208.410 48.170 208.580 ;
        RECT 45.235 207.930 45.700 208.240 ;
        RECT 45.880 207.930 46.405 208.240 ;
        RECT 44.765 207.550 45.995 207.750 ;
        RECT 44.835 207.000 45.505 207.370 ;
        RECT 45.685 207.180 45.995 207.550 ;
        RECT 46.175 207.290 46.405 207.930 ;
        RECT 46.585 207.910 46.885 208.240 ;
        RECT 46.585 207.000 46.875 207.730 ;
        RECT 47.065 207.675 47.235 208.410 ;
        RECT 47.510 208.240 47.680 208.410 ;
        RECT 48.430 208.240 48.675 208.530 ;
        RECT 48.845 208.410 49.175 208.700 ;
        RECT 49.435 208.240 49.605 208.800 ;
        RECT 49.855 208.410 50.115 209.550 ;
        RECT 50.375 208.620 50.545 209.380 ;
        RECT 50.760 208.790 51.090 209.550 ;
        RECT 50.375 208.450 51.090 208.620 ;
        RECT 51.260 208.475 51.515 209.380 ;
        RECT 47.405 207.910 47.680 208.240 ;
        RECT 47.850 207.910 48.675 208.240 ;
        RECT 48.890 207.910 49.605 208.240 ;
        RECT 49.775 207.990 50.110 208.240 ;
        RECT 47.510 207.740 47.680 207.910 ;
        RECT 49.355 207.820 49.605 207.910 ;
        RECT 50.285 207.900 50.640 208.270 ;
        RECT 50.920 208.240 51.090 208.450 ;
        RECT 50.920 207.910 51.175 208.240 ;
        RECT 47.065 207.330 47.340 207.675 ;
        RECT 47.510 207.570 49.175 207.740 ;
        RECT 47.530 207.000 47.905 207.400 ;
        RECT 48.075 207.220 48.245 207.570 ;
        RECT 48.415 207.000 48.745 207.400 ;
        RECT 48.915 207.170 49.175 207.570 ;
        RECT 49.355 207.400 49.685 207.820 ;
        RECT 49.855 207.000 50.115 207.820 ;
        RECT 50.920 207.720 51.090 207.910 ;
        RECT 51.345 207.745 51.515 208.475 ;
        RECT 51.690 208.400 51.950 209.550 ;
        RECT 52.585 208.385 52.875 209.550 ;
        RECT 53.045 208.960 53.745 209.380 ;
        RECT 53.945 209.190 54.275 209.550 ;
        RECT 54.445 208.960 54.775 209.360 ;
        RECT 53.045 208.730 54.775 208.960 ;
        RECT 50.375 207.550 51.090 207.720 ;
        RECT 50.375 207.170 50.545 207.550 ;
        RECT 50.760 207.000 51.090 207.380 ;
        RECT 51.260 207.170 51.515 207.745 ;
        RECT 51.690 207.000 51.950 207.840 ;
        RECT 53.045 207.760 53.250 208.730 ;
        RECT 53.420 207.990 53.750 208.530 ;
        RECT 53.925 208.240 54.250 208.530 ;
        RECT 54.445 208.510 54.775 208.730 ;
        RECT 54.945 208.240 55.115 209.210 ;
        RECT 55.295 208.490 55.625 209.550 ;
        RECT 55.805 208.830 56.265 209.380 ;
        RECT 56.455 208.830 56.785 209.550 ;
        RECT 53.925 207.910 54.420 208.240 ;
        RECT 54.740 207.910 55.115 208.240 ;
        RECT 55.325 207.910 55.635 208.240 ;
        RECT 52.585 207.000 52.875 207.725 ;
        RECT 53.045 207.170 53.755 207.760 ;
        RECT 54.265 207.530 55.625 207.740 ;
        RECT 54.265 207.170 54.595 207.530 ;
        RECT 54.795 207.000 55.125 207.360 ;
        RECT 55.295 207.170 55.625 207.530 ;
        RECT 55.805 207.460 56.055 208.830 ;
        RECT 56.985 208.660 57.285 209.210 ;
        RECT 57.455 208.880 57.735 209.550 ;
        RECT 56.345 208.490 57.285 208.660 ;
        RECT 56.345 208.240 56.515 208.490 ;
        RECT 57.655 208.240 57.920 208.600 ;
        RECT 59.075 208.410 59.325 209.550 ;
        RECT 56.225 207.910 56.515 208.240 ;
        RECT 56.685 207.990 57.025 208.240 ;
        RECT 57.245 207.990 57.920 208.240 ;
        RECT 59.495 208.360 59.745 209.240 ;
        RECT 59.915 208.410 60.220 209.550 ;
        RECT 60.560 209.170 60.890 209.550 ;
        RECT 61.070 209.000 61.240 209.290 ;
        RECT 61.410 209.090 61.660 209.550 ;
        RECT 60.440 208.830 61.240 209.000 ;
        RECT 61.830 209.040 62.700 209.380 ;
        RECT 56.345 207.820 56.515 207.910 ;
        RECT 56.345 207.630 57.735 207.820 ;
        RECT 55.805 207.170 56.365 207.460 ;
        RECT 56.535 207.000 56.785 207.460 ;
        RECT 57.405 207.270 57.735 207.630 ;
        RECT 59.075 207.000 59.325 207.755 ;
        RECT 59.495 207.710 59.700 208.360 ;
        RECT 60.440 208.240 60.610 208.830 ;
        RECT 61.830 208.660 62.000 209.040 ;
        RECT 62.935 208.920 63.105 209.380 ;
        RECT 63.275 209.090 63.645 209.550 ;
        RECT 63.940 208.950 64.110 209.290 ;
        RECT 64.280 209.120 64.610 209.550 ;
        RECT 64.845 208.950 65.015 209.290 ;
        RECT 60.780 208.490 62.000 208.660 ;
        RECT 62.170 208.580 62.630 208.870 ;
        RECT 62.935 208.750 63.495 208.920 ;
        RECT 63.940 208.780 65.015 208.950 ;
        RECT 65.185 209.050 65.865 209.380 ;
        RECT 66.080 209.050 66.330 209.380 ;
        RECT 66.500 209.090 66.750 209.550 ;
        RECT 63.325 208.610 63.495 208.750 ;
        RECT 62.170 208.570 63.135 208.580 ;
        RECT 61.830 208.400 62.000 208.490 ;
        RECT 62.460 208.410 63.135 208.570 ;
        RECT 59.870 208.210 60.610 208.240 ;
        RECT 59.870 207.910 60.785 208.210 ;
        RECT 60.460 207.735 60.785 207.910 ;
        RECT 59.495 207.180 59.745 207.710 ;
        RECT 59.915 207.000 60.220 207.460 ;
        RECT 60.465 207.380 60.785 207.735 ;
        RECT 60.955 207.950 61.495 208.320 ;
        RECT 61.830 208.230 62.235 208.400 ;
        RECT 60.955 207.550 61.195 207.950 ;
        RECT 61.675 207.780 61.895 208.060 ;
        RECT 61.365 207.610 61.895 207.780 ;
        RECT 61.365 207.380 61.535 207.610 ;
        RECT 62.065 207.450 62.235 208.230 ;
        RECT 62.405 207.620 62.755 208.240 ;
        RECT 62.925 207.620 63.135 208.410 ;
        RECT 63.325 208.440 64.825 208.610 ;
        RECT 63.325 207.750 63.495 208.440 ;
        RECT 65.185 208.270 65.355 209.050 ;
        RECT 66.160 208.920 66.330 209.050 ;
        RECT 63.665 208.100 65.355 208.270 ;
        RECT 65.525 208.490 65.990 208.880 ;
        RECT 66.160 208.750 66.555 208.920 ;
        RECT 63.665 207.920 63.835 208.100 ;
        RECT 60.465 207.210 61.535 207.380 ;
        RECT 61.705 207.000 61.895 207.440 ;
        RECT 62.065 207.170 63.015 207.450 ;
        RECT 63.325 207.360 63.585 207.750 ;
        RECT 64.005 207.680 64.795 207.930 ;
        RECT 63.235 207.190 63.585 207.360 ;
        RECT 63.795 207.000 64.125 207.460 ;
        RECT 65.000 207.390 65.170 208.100 ;
        RECT 65.525 207.900 65.695 208.490 ;
        RECT 65.340 207.680 65.695 207.900 ;
        RECT 65.865 207.680 66.215 208.300 ;
        RECT 66.385 207.390 66.555 208.750 ;
        RECT 66.920 208.580 67.245 209.365 ;
        RECT 66.725 207.530 67.185 208.580 ;
        RECT 65.000 207.220 65.855 207.390 ;
        RECT 66.060 207.220 66.555 207.390 ;
        RECT 66.725 207.000 67.055 207.360 ;
        RECT 67.415 207.260 67.585 209.380 ;
        RECT 67.755 209.050 68.085 209.550 ;
        RECT 68.255 208.880 68.510 209.380 ;
        RECT 67.760 208.710 68.510 208.880 ;
        RECT 69.605 208.960 70.305 209.380 ;
        RECT 70.505 209.190 70.835 209.550 ;
        RECT 71.005 208.960 71.335 209.360 ;
        RECT 69.605 208.730 71.335 208.960 ;
        RECT 67.760 207.720 67.990 208.710 ;
        RECT 68.160 207.890 68.510 208.540 ;
        RECT 69.605 207.760 69.810 208.730 ;
        RECT 69.980 207.990 70.310 208.530 ;
        RECT 70.485 208.240 70.810 208.530 ;
        RECT 71.005 208.510 71.335 208.730 ;
        RECT 71.505 208.240 71.675 209.165 ;
        RECT 71.855 208.490 72.185 209.550 ;
        RECT 72.375 208.490 72.705 209.340 ;
        RECT 70.485 207.910 70.980 208.240 ;
        RECT 71.300 207.910 71.675 208.240 ;
        RECT 71.885 207.910 72.195 208.240 ;
        RECT 67.760 207.550 68.510 207.720 ;
        RECT 67.755 207.000 68.085 207.380 ;
        RECT 68.255 207.260 68.510 207.550 ;
        RECT 69.605 207.170 70.315 207.760 ;
        RECT 70.825 207.530 72.185 207.740 ;
        RECT 70.825 207.170 71.155 207.530 ;
        RECT 71.355 207.000 71.685 207.360 ;
        RECT 71.855 207.170 72.185 207.530 ;
        RECT 72.375 207.725 72.565 208.490 ;
        RECT 72.875 208.410 73.125 209.550 ;
        RECT 73.315 208.910 73.565 209.330 ;
        RECT 73.795 209.080 74.125 209.550 ;
        RECT 74.355 208.910 74.605 209.330 ;
        RECT 73.315 208.740 74.605 208.910 ;
        RECT 74.785 208.910 75.115 209.340 ;
        RECT 74.785 208.740 75.240 208.910 ;
        RECT 73.305 208.240 73.520 208.570 ;
        RECT 72.735 207.910 73.045 208.240 ;
        RECT 73.215 207.910 73.520 208.240 ;
        RECT 73.695 207.910 73.980 208.570 ;
        RECT 74.175 207.910 74.440 208.570 ;
        RECT 74.655 207.910 74.900 208.570 ;
        RECT 72.875 207.740 73.045 207.910 ;
        RECT 75.070 207.740 75.240 208.740 ;
        RECT 75.590 208.410 75.910 209.550 ;
        RECT 76.090 208.240 76.285 209.290 ;
        RECT 76.465 208.700 76.795 209.380 ;
        RECT 76.995 208.750 77.250 209.550 ;
        RECT 76.465 208.420 76.815 208.700 ;
        RECT 75.650 208.190 75.910 208.240 ;
        RECT 75.645 208.020 75.910 208.190 ;
        RECT 75.650 207.910 75.910 208.020 ;
        RECT 76.090 207.910 76.475 208.240 ;
        RECT 76.645 208.040 76.815 208.420 ;
        RECT 77.005 208.210 77.250 208.570 ;
        RECT 78.345 208.385 78.635 209.550 ;
        RECT 79.730 208.830 80.065 209.340 ;
        RECT 76.645 207.870 77.165 208.040 ;
        RECT 72.375 207.215 72.705 207.725 ;
        RECT 72.875 207.570 75.240 207.740 ;
        RECT 72.875 207.000 73.205 207.400 ;
        RECT 74.255 207.230 74.585 207.570 ;
        RECT 75.590 207.530 76.805 207.700 ;
        RECT 74.755 207.000 75.085 207.400 ;
        RECT 75.590 207.180 75.880 207.530 ;
        RECT 76.075 207.000 76.405 207.360 ;
        RECT 76.575 207.225 76.805 207.530 ;
        RECT 76.995 207.305 77.165 207.870 ;
        RECT 78.345 207.000 78.635 207.725 ;
        RECT 79.730 207.475 79.985 208.830 ;
        RECT 80.315 208.750 80.645 209.550 ;
        RECT 80.890 208.960 81.175 209.380 ;
        RECT 81.430 209.130 81.760 209.550 ;
        RECT 81.985 209.210 83.145 209.380 ;
        RECT 81.985 208.960 82.315 209.210 ;
        RECT 80.890 208.790 82.315 208.960 ;
        RECT 82.545 208.580 82.715 209.040 ;
        RECT 82.975 208.710 83.145 209.210 ;
        RECT 84.325 208.960 85.025 209.380 ;
        RECT 85.225 209.190 85.555 209.550 ;
        RECT 85.725 208.960 86.055 209.360 ;
        RECT 84.325 208.730 86.055 208.960 ;
        RECT 80.345 208.410 82.715 208.580 ;
        RECT 80.345 208.240 80.515 208.410 ;
        RECT 82.965 208.360 83.175 208.530 ;
        RECT 82.965 208.240 83.170 208.360 ;
        RECT 80.210 207.910 80.515 208.240 ;
        RECT 80.710 208.190 80.960 208.240 ;
        RECT 81.170 208.190 81.440 208.240 ;
        RECT 80.705 208.020 80.960 208.190 ;
        RECT 81.165 208.020 81.440 208.190 ;
        RECT 80.710 207.910 80.960 208.020 ;
        RECT 80.345 207.740 80.515 207.910 ;
        RECT 80.345 207.570 80.905 207.740 ;
        RECT 81.170 207.580 81.440 208.020 ;
        RECT 81.630 207.850 81.920 208.240 ;
        RECT 81.625 207.680 81.920 207.850 ;
        RECT 81.630 207.580 81.920 207.680 ;
        RECT 82.090 207.575 82.510 208.240 ;
        RECT 82.820 207.910 83.170 208.240 ;
        RECT 84.325 207.760 84.530 208.730 ;
        RECT 84.700 207.990 85.030 208.530 ;
        RECT 85.205 208.240 85.530 208.530 ;
        RECT 85.725 208.510 86.055 208.730 ;
        RECT 86.225 208.240 86.395 209.165 ;
        RECT 86.575 208.490 86.905 209.550 ;
        RECT 87.090 208.830 87.425 209.340 ;
        RECT 85.205 207.910 85.700 208.240 ;
        RECT 86.020 207.910 86.395 208.240 ;
        RECT 86.605 207.910 86.915 208.240 ;
        RECT 79.730 207.215 80.065 207.475 ;
        RECT 80.735 207.400 80.905 207.570 ;
        RECT 80.235 207.000 80.565 207.400 ;
        RECT 80.735 207.230 82.350 207.400 ;
        RECT 82.895 207.000 83.225 207.720 ;
        RECT 84.325 207.170 85.035 207.760 ;
        RECT 85.545 207.530 86.905 207.740 ;
        RECT 85.545 207.170 85.875 207.530 ;
        RECT 86.075 207.000 86.405 207.360 ;
        RECT 86.575 207.170 86.905 207.530 ;
        RECT 87.090 207.475 87.345 208.830 ;
        RECT 87.675 208.750 88.005 209.550 ;
        RECT 88.250 208.960 88.535 209.380 ;
        RECT 88.790 209.130 89.120 209.550 ;
        RECT 89.345 209.210 90.505 209.380 ;
        RECT 89.345 208.960 89.675 209.210 ;
        RECT 88.250 208.790 89.675 208.960 ;
        RECT 89.905 208.580 90.075 209.040 ;
        RECT 90.335 208.710 90.505 209.210 ;
        RECT 87.705 208.410 90.075 208.580 ;
        RECT 87.705 208.240 87.875 208.410 ;
        RECT 90.325 208.240 90.530 208.530 ;
        RECT 87.570 207.910 87.875 208.240 ;
        RECT 88.070 208.190 88.320 208.240 ;
        RECT 88.530 208.190 88.800 208.240 ;
        RECT 88.990 208.190 89.280 208.240 ;
        RECT 88.065 208.020 88.320 208.190 ;
        RECT 88.525 208.020 88.800 208.190 ;
        RECT 88.985 208.020 89.280 208.190 ;
        RECT 88.070 207.910 88.320 208.020 ;
        RECT 87.705 207.740 87.875 207.910 ;
        RECT 87.705 207.570 88.265 207.740 ;
        RECT 88.530 207.580 88.800 208.020 ;
        RECT 88.990 207.580 89.280 208.020 ;
        RECT 89.450 207.575 89.870 208.240 ;
        RECT 90.180 208.190 90.530 208.240 ;
        RECT 91.685 208.410 91.945 209.380 ;
        RECT 92.140 209.140 92.470 209.550 ;
        RECT 92.670 208.960 92.840 209.380 ;
        RECT 93.055 209.140 93.725 209.550 ;
        RECT 93.960 208.960 94.130 209.380 ;
        RECT 94.435 209.110 94.765 209.550 ;
        RECT 92.115 208.790 94.130 208.960 ;
        RECT 94.935 208.930 95.110 209.380 ;
        RECT 90.180 208.020 90.535 208.190 ;
        RECT 90.180 207.910 90.530 208.020 ;
        RECT 91.685 207.720 91.855 208.410 ;
        RECT 92.115 208.240 92.285 208.790 ;
        RECT 92.025 207.910 92.285 208.240 ;
        RECT 87.090 207.215 87.425 207.475 ;
        RECT 88.095 207.400 88.265 207.570 ;
        RECT 87.595 207.000 87.925 207.400 ;
        RECT 88.095 207.230 89.710 207.400 ;
        RECT 90.255 207.000 90.585 207.720 ;
        RECT 91.685 207.255 92.025 207.720 ;
        RECT 92.455 207.580 92.795 208.610 ;
        RECT 92.985 207.850 93.255 208.610 ;
        RECT 92.985 207.680 93.295 207.850 ;
        RECT 91.690 207.210 92.025 207.255 ;
        RECT 92.195 207.000 92.525 207.380 ;
        RECT 92.985 207.335 93.255 207.680 ;
        RECT 93.480 207.335 93.760 208.610 ;
        RECT 93.960 207.500 94.130 208.790 ;
        RECT 94.480 208.760 95.110 208.930 ;
        RECT 94.480 208.240 94.650 208.760 ;
        RECT 94.300 207.910 94.650 208.240 ;
        RECT 94.830 207.910 95.195 208.590 ;
        RECT 95.365 208.410 95.625 209.380 ;
        RECT 95.820 209.140 96.150 209.550 ;
        RECT 96.350 208.960 96.520 209.380 ;
        RECT 96.735 209.140 97.405 209.550 ;
        RECT 97.640 208.960 97.810 209.380 ;
        RECT 98.115 209.110 98.445 209.550 ;
        RECT 95.795 208.790 97.810 208.960 ;
        RECT 98.615 208.930 98.790 209.380 ;
        RECT 94.480 207.740 94.650 207.910 ;
        RECT 94.480 207.570 95.110 207.740 ;
        RECT 93.960 207.170 94.190 207.500 ;
        RECT 94.435 207.000 94.765 207.380 ;
        RECT 94.935 207.170 95.110 207.570 ;
        RECT 95.365 207.720 95.535 208.410 ;
        RECT 95.795 208.240 95.965 208.790 ;
        RECT 95.705 207.910 95.965 208.240 ;
        RECT 95.365 207.255 95.705 207.720 ;
        RECT 96.135 207.580 96.475 208.610 ;
        RECT 96.665 207.510 96.935 208.610 ;
        RECT 95.370 207.210 95.705 207.255 ;
        RECT 95.875 207.000 96.205 207.380 ;
        RECT 96.665 207.340 96.975 207.510 ;
        RECT 96.665 207.335 96.935 207.340 ;
        RECT 97.160 207.335 97.440 208.610 ;
        RECT 97.640 207.500 97.810 208.790 ;
        RECT 98.160 208.760 98.790 208.930 ;
        RECT 98.160 208.240 98.330 208.760 ;
        RECT 97.980 207.910 98.330 208.240 ;
        RECT 98.510 207.910 98.875 208.590 ;
        RECT 99.055 208.490 99.385 209.340 ;
        RECT 98.160 207.740 98.330 207.910 ;
        RECT 98.160 207.570 98.790 207.740 ;
        RECT 97.640 207.170 97.870 207.500 ;
        RECT 98.115 207.000 98.445 207.380 ;
        RECT 98.615 207.170 98.790 207.570 ;
        RECT 99.055 207.725 99.245 208.490 ;
        RECT 99.555 208.410 99.805 209.550 ;
        RECT 99.995 208.910 100.245 209.330 ;
        RECT 100.475 209.080 100.805 209.550 ;
        RECT 101.035 208.910 101.285 209.330 ;
        RECT 99.995 208.740 101.285 208.910 ;
        RECT 101.465 208.910 101.795 209.340 ;
        RECT 101.465 208.740 101.920 208.910 ;
        RECT 99.985 208.240 100.200 208.570 ;
        RECT 99.415 207.910 99.725 208.240 ;
        RECT 99.895 207.910 100.200 208.240 ;
        RECT 100.375 207.910 100.660 208.570 ;
        RECT 100.855 207.910 101.120 208.570 ;
        RECT 101.335 207.910 101.580 208.570 ;
        RECT 99.555 207.740 99.725 207.910 ;
        RECT 101.750 207.740 101.920 208.740 ;
        RECT 99.055 207.215 99.385 207.725 ;
        RECT 99.555 207.570 101.920 207.740 ;
        RECT 102.265 208.580 102.535 209.350 ;
        RECT 102.705 208.770 103.035 209.550 ;
        RECT 103.240 208.945 103.425 209.350 ;
        RECT 103.595 209.125 103.930 209.550 ;
        RECT 103.240 208.770 103.905 208.945 ;
        RECT 102.265 208.410 103.395 208.580 ;
        RECT 99.555 207.000 99.885 207.400 ;
        RECT 100.935 207.230 101.265 207.570 ;
        RECT 102.265 207.500 102.435 208.410 ;
        RECT 102.605 207.660 102.965 208.240 ;
        RECT 103.145 207.910 103.395 208.410 ;
        RECT 103.565 207.740 103.905 208.770 ;
        RECT 104.105 208.385 104.395 209.550 ;
        RECT 104.565 208.410 104.825 209.550 ;
        RECT 105.065 209.040 106.680 209.370 ;
        RECT 105.075 208.240 105.245 208.800 ;
        RECT 105.505 208.700 106.680 208.870 ;
        RECT 106.850 208.750 107.130 209.550 ;
        RECT 105.505 208.410 105.835 208.700 ;
        RECT 106.510 208.580 106.680 208.700 ;
        RECT 106.005 208.240 106.250 208.530 ;
        RECT 106.510 208.410 107.170 208.580 ;
        RECT 107.340 208.410 107.615 209.380 ;
        RECT 107.790 208.880 108.045 209.380 ;
        RECT 108.215 209.050 108.545 209.550 ;
        RECT 107.790 208.710 108.540 208.880 ;
        RECT 107.000 208.240 107.170 208.410 ;
        RECT 104.570 207.990 104.905 208.240 ;
        RECT 105.075 207.910 105.790 208.240 ;
        RECT 106.005 207.910 106.830 208.240 ;
        RECT 107.000 207.910 107.275 208.240 ;
        RECT 105.075 207.820 105.325 207.910 ;
        RECT 103.220 207.570 103.905 207.740 ;
        RECT 101.435 207.000 101.765 207.400 ;
        RECT 102.265 207.170 102.525 207.500 ;
        RECT 102.735 207.000 103.010 207.480 ;
        RECT 103.220 207.170 103.425 207.570 ;
        RECT 103.595 207.000 103.930 207.400 ;
        RECT 104.105 207.000 104.395 207.725 ;
        RECT 104.565 207.000 104.825 207.820 ;
        RECT 104.995 207.400 105.325 207.820 ;
        RECT 107.000 207.740 107.170 207.910 ;
        RECT 105.505 207.570 107.170 207.740 ;
        RECT 107.445 207.675 107.615 208.410 ;
        RECT 107.790 207.890 108.140 208.540 ;
        RECT 108.310 207.720 108.540 208.710 ;
        RECT 105.505 207.170 105.765 207.570 ;
        RECT 105.935 207.000 106.265 207.400 ;
        RECT 106.435 207.220 106.605 207.570 ;
        RECT 106.775 207.000 107.150 207.400 ;
        RECT 107.340 207.330 107.615 207.675 ;
        RECT 107.790 207.550 108.540 207.720 ;
        RECT 107.790 207.260 108.045 207.550 ;
        RECT 108.215 207.000 108.545 207.380 ;
        RECT 108.715 207.260 108.885 209.380 ;
        RECT 109.055 208.580 109.380 209.365 ;
        RECT 109.550 209.090 109.800 209.550 ;
        RECT 109.970 209.050 110.220 209.380 ;
        RECT 110.435 209.050 111.115 209.380 ;
        RECT 109.970 208.920 110.140 209.050 ;
        RECT 109.745 208.750 110.140 208.920 ;
        RECT 109.115 207.530 109.575 208.580 ;
        RECT 109.745 207.390 109.915 208.750 ;
        RECT 110.310 208.490 110.775 208.880 ;
        RECT 110.085 207.680 110.435 208.300 ;
        RECT 110.605 207.900 110.775 208.490 ;
        RECT 110.945 208.270 111.115 209.050 ;
        RECT 111.285 208.950 111.455 209.290 ;
        RECT 111.690 209.120 112.020 209.550 ;
        RECT 112.190 208.950 112.360 209.290 ;
        RECT 112.655 209.090 113.025 209.550 ;
        RECT 111.285 208.780 112.360 208.950 ;
        RECT 113.195 208.920 113.365 209.380 ;
        RECT 113.600 209.040 114.470 209.380 ;
        RECT 114.640 209.090 114.890 209.550 ;
        RECT 112.805 208.750 113.365 208.920 ;
        RECT 112.805 208.610 112.975 208.750 ;
        RECT 111.475 208.440 112.975 208.610 ;
        RECT 113.670 208.580 114.130 208.870 ;
        RECT 110.945 208.100 112.635 208.270 ;
        RECT 110.605 207.680 110.960 207.900 ;
        RECT 111.130 207.390 111.300 208.100 ;
        RECT 111.505 207.680 112.295 207.930 ;
        RECT 112.465 207.920 112.635 208.100 ;
        RECT 112.805 207.750 112.975 208.440 ;
        RECT 109.245 207.000 109.575 207.360 ;
        RECT 109.745 207.220 110.240 207.390 ;
        RECT 110.445 207.220 111.300 207.390 ;
        RECT 112.175 207.000 112.505 207.460 ;
        RECT 112.715 207.360 112.975 207.750 ;
        RECT 113.165 208.570 114.130 208.580 ;
        RECT 114.300 208.660 114.470 209.040 ;
        RECT 115.060 209.000 115.230 209.290 ;
        RECT 115.410 209.170 115.740 209.550 ;
        RECT 115.060 208.830 115.860 209.000 ;
        RECT 113.165 208.410 113.840 208.570 ;
        RECT 114.300 208.490 115.520 208.660 ;
        RECT 113.165 207.620 113.375 208.410 ;
        RECT 114.300 208.400 114.470 208.490 ;
        RECT 113.545 207.620 113.895 208.240 ;
        RECT 114.065 208.230 114.470 208.400 ;
        RECT 114.065 207.450 114.235 208.230 ;
        RECT 114.405 207.780 114.625 208.060 ;
        RECT 114.805 207.950 115.345 208.320 ;
        RECT 115.690 208.240 115.860 208.830 ;
        RECT 116.080 208.410 116.385 209.550 ;
        RECT 116.555 208.360 116.810 209.240 ;
        RECT 117.190 208.580 117.520 209.380 ;
        RECT 117.690 208.750 118.020 209.550 ;
        RECT 118.320 208.580 118.650 209.380 ;
        RECT 119.295 208.750 119.545 209.550 ;
        RECT 117.190 208.410 119.625 208.580 ;
        RECT 119.815 208.410 119.985 209.550 ;
        RECT 120.155 208.410 120.495 209.380 ;
        RECT 120.670 208.880 120.925 209.380 ;
        RECT 121.095 209.050 121.425 209.550 ;
        RECT 120.670 208.710 121.420 208.880 ;
        RECT 115.690 208.210 116.430 208.240 ;
        RECT 114.405 207.610 114.935 207.780 ;
        RECT 112.715 207.190 113.065 207.360 ;
        RECT 113.285 207.170 114.235 207.450 ;
        RECT 114.405 207.000 114.595 207.440 ;
        RECT 114.765 207.380 114.935 207.610 ;
        RECT 115.105 207.550 115.345 207.950 ;
        RECT 115.515 207.910 116.430 208.210 ;
        RECT 115.515 207.735 115.840 207.910 ;
        RECT 115.515 207.380 115.835 207.735 ;
        RECT 116.600 207.710 116.810 208.360 ;
        RECT 116.985 207.990 117.335 208.240 ;
        RECT 117.520 207.780 117.690 208.410 ;
        RECT 117.860 207.990 118.190 208.190 ;
        RECT 118.360 207.990 118.690 208.190 ;
        RECT 118.860 207.990 119.280 208.190 ;
        RECT 119.455 208.160 119.625 208.410 ;
        RECT 119.455 207.990 120.150 208.160 ;
        RECT 114.765 207.210 115.835 207.380 ;
        RECT 116.080 207.000 116.385 207.460 ;
        RECT 116.555 207.180 116.810 207.710 ;
        RECT 117.190 207.170 117.690 207.780 ;
        RECT 118.320 207.650 119.545 207.820 ;
        RECT 120.320 207.800 120.495 208.410 ;
        RECT 120.670 207.890 121.020 208.540 ;
        RECT 118.320 207.170 118.650 207.650 ;
        RECT 118.820 207.000 119.045 207.460 ;
        RECT 119.215 207.170 119.545 207.650 ;
        RECT 119.735 207.000 119.985 207.800 ;
        RECT 120.155 207.170 120.495 207.800 ;
        RECT 121.190 207.720 121.420 208.710 ;
        RECT 120.670 207.550 121.420 207.720 ;
        RECT 120.670 207.260 120.925 207.550 ;
        RECT 121.095 207.000 121.425 207.380 ;
        RECT 121.595 207.260 121.765 209.380 ;
        RECT 121.935 208.580 122.260 209.365 ;
        RECT 122.430 209.090 122.680 209.550 ;
        RECT 122.850 209.050 123.100 209.380 ;
        RECT 123.315 209.050 123.995 209.380 ;
        RECT 122.850 208.920 123.020 209.050 ;
        RECT 122.625 208.750 123.020 208.920 ;
        RECT 121.995 207.530 122.455 208.580 ;
        RECT 122.625 207.390 122.795 208.750 ;
        RECT 123.190 208.490 123.655 208.880 ;
        RECT 122.965 207.680 123.315 208.300 ;
        RECT 123.485 207.900 123.655 208.490 ;
        RECT 123.825 208.270 123.995 209.050 ;
        RECT 124.165 208.950 124.335 209.290 ;
        RECT 124.570 209.120 124.900 209.550 ;
        RECT 125.070 208.950 125.240 209.290 ;
        RECT 125.535 209.090 125.905 209.550 ;
        RECT 124.165 208.780 125.240 208.950 ;
        RECT 126.075 208.920 126.245 209.380 ;
        RECT 126.480 209.040 127.350 209.380 ;
        RECT 127.520 209.090 127.770 209.550 ;
        RECT 125.685 208.750 126.245 208.920 ;
        RECT 125.685 208.610 125.855 208.750 ;
        RECT 124.355 208.440 125.855 208.610 ;
        RECT 126.550 208.580 127.010 208.870 ;
        RECT 123.825 208.100 125.515 208.270 ;
        RECT 123.485 207.680 123.840 207.900 ;
        RECT 124.010 207.390 124.180 208.100 ;
        RECT 124.385 207.680 125.175 207.930 ;
        RECT 125.345 207.920 125.515 208.100 ;
        RECT 125.685 207.750 125.855 208.440 ;
        RECT 122.125 207.000 122.455 207.360 ;
        RECT 122.625 207.220 123.120 207.390 ;
        RECT 123.325 207.220 124.180 207.390 ;
        RECT 125.055 207.000 125.385 207.460 ;
        RECT 125.595 207.360 125.855 207.750 ;
        RECT 126.045 208.570 127.010 208.580 ;
        RECT 127.180 208.660 127.350 209.040 ;
        RECT 127.940 209.000 128.110 209.290 ;
        RECT 128.290 209.170 128.620 209.550 ;
        RECT 127.940 208.830 128.740 209.000 ;
        RECT 126.045 208.410 126.720 208.570 ;
        RECT 127.180 208.490 128.400 208.660 ;
        RECT 126.045 207.620 126.255 208.410 ;
        RECT 127.180 208.400 127.350 208.490 ;
        RECT 126.425 207.620 126.775 208.240 ;
        RECT 126.945 208.230 127.350 208.400 ;
        RECT 126.945 207.450 127.115 208.230 ;
        RECT 127.285 207.780 127.505 208.060 ;
        RECT 127.685 207.950 128.225 208.320 ;
        RECT 128.570 208.240 128.740 208.830 ;
        RECT 128.960 208.410 129.265 209.550 ;
        RECT 129.435 208.360 129.690 209.240 ;
        RECT 129.865 208.385 130.155 209.550 ;
        RECT 130.330 208.880 130.585 209.380 ;
        RECT 130.755 209.050 131.085 209.550 ;
        RECT 130.330 208.710 131.080 208.880 ;
        RECT 128.570 208.210 129.310 208.240 ;
        RECT 127.285 207.610 127.815 207.780 ;
        RECT 125.595 207.190 125.945 207.360 ;
        RECT 126.165 207.170 127.115 207.450 ;
        RECT 127.285 207.000 127.475 207.440 ;
        RECT 127.645 207.380 127.815 207.610 ;
        RECT 127.985 207.550 128.225 207.950 ;
        RECT 128.395 207.910 129.310 208.210 ;
        RECT 128.395 207.735 128.720 207.910 ;
        RECT 128.395 207.380 128.715 207.735 ;
        RECT 129.480 207.710 129.690 208.360 ;
        RECT 130.330 207.890 130.680 208.540 ;
        RECT 127.645 207.210 128.715 207.380 ;
        RECT 128.960 207.000 129.265 207.460 ;
        RECT 129.435 207.180 129.690 207.710 ;
        RECT 129.865 207.000 130.155 207.725 ;
        RECT 130.850 207.720 131.080 208.710 ;
        RECT 130.330 207.550 131.080 207.720 ;
        RECT 130.330 207.260 130.585 207.550 ;
        RECT 130.755 207.000 131.085 207.380 ;
        RECT 131.255 207.260 131.425 209.380 ;
        RECT 131.595 208.580 131.920 209.365 ;
        RECT 132.090 209.090 132.340 209.550 ;
        RECT 132.510 209.050 132.760 209.380 ;
        RECT 132.975 209.050 133.655 209.380 ;
        RECT 132.510 208.920 132.680 209.050 ;
        RECT 132.285 208.750 132.680 208.920 ;
        RECT 131.655 207.530 132.115 208.580 ;
        RECT 132.285 207.390 132.455 208.750 ;
        RECT 132.850 208.490 133.315 208.880 ;
        RECT 132.625 207.680 132.975 208.300 ;
        RECT 133.145 207.900 133.315 208.490 ;
        RECT 133.485 208.270 133.655 209.050 ;
        RECT 133.825 208.950 133.995 209.290 ;
        RECT 134.230 209.120 134.560 209.550 ;
        RECT 134.730 208.950 134.900 209.290 ;
        RECT 135.195 209.090 135.565 209.550 ;
        RECT 133.825 208.780 134.900 208.950 ;
        RECT 135.735 208.920 135.905 209.380 ;
        RECT 136.140 209.040 137.010 209.380 ;
        RECT 137.180 209.090 137.430 209.550 ;
        RECT 135.345 208.750 135.905 208.920 ;
        RECT 135.345 208.610 135.515 208.750 ;
        RECT 134.015 208.440 135.515 208.610 ;
        RECT 136.210 208.580 136.670 208.870 ;
        RECT 133.485 208.100 135.175 208.270 ;
        RECT 133.145 207.680 133.500 207.900 ;
        RECT 133.670 207.390 133.840 208.100 ;
        RECT 134.045 207.680 134.835 207.930 ;
        RECT 135.005 207.920 135.175 208.100 ;
        RECT 135.345 207.750 135.515 208.440 ;
        RECT 131.785 207.000 132.115 207.360 ;
        RECT 132.285 207.220 132.780 207.390 ;
        RECT 132.985 207.220 133.840 207.390 ;
        RECT 134.715 207.000 135.045 207.460 ;
        RECT 135.255 207.360 135.515 207.750 ;
        RECT 135.705 208.570 136.670 208.580 ;
        RECT 136.840 208.660 137.010 209.040 ;
        RECT 137.600 209.000 137.770 209.290 ;
        RECT 137.950 209.170 138.280 209.550 ;
        RECT 137.600 208.830 138.400 209.000 ;
        RECT 135.705 208.410 136.380 208.570 ;
        RECT 136.840 208.490 138.060 208.660 ;
        RECT 135.705 207.620 135.915 208.410 ;
        RECT 136.840 208.400 137.010 208.490 ;
        RECT 136.085 207.620 136.435 208.240 ;
        RECT 136.605 208.230 137.010 208.400 ;
        RECT 136.605 207.450 136.775 208.230 ;
        RECT 136.945 207.780 137.165 208.060 ;
        RECT 137.345 207.950 137.885 208.320 ;
        RECT 138.230 208.240 138.400 208.830 ;
        RECT 138.620 208.410 138.925 209.550 ;
        RECT 139.095 208.360 139.350 209.240 ;
        RECT 139.525 208.460 140.735 209.550 ;
        RECT 138.230 208.210 138.970 208.240 ;
        RECT 136.945 207.610 137.475 207.780 ;
        RECT 135.255 207.190 135.605 207.360 ;
        RECT 135.825 207.170 136.775 207.450 ;
        RECT 136.945 207.000 137.135 207.440 ;
        RECT 137.305 207.380 137.475 207.610 ;
        RECT 137.645 207.550 137.885 207.950 ;
        RECT 138.055 207.910 138.970 208.210 ;
        RECT 138.055 207.735 138.380 207.910 ;
        RECT 138.055 207.380 138.375 207.735 ;
        RECT 139.140 207.710 139.350 208.360 ;
        RECT 137.305 207.210 138.375 207.380 ;
        RECT 138.620 207.000 138.925 207.460 ;
        RECT 139.095 207.180 139.350 207.710 ;
        RECT 139.525 207.750 140.045 208.290 ;
        RECT 140.215 207.920 140.735 208.460 ;
        RECT 140.995 208.620 141.165 209.380 ;
        RECT 141.380 208.790 141.710 209.550 ;
        RECT 140.995 208.450 141.710 208.620 ;
        RECT 141.880 208.475 142.135 209.380 ;
        RECT 140.905 207.900 141.260 208.270 ;
        RECT 141.540 208.240 141.710 208.450 ;
        RECT 141.540 207.910 141.795 208.240 ;
        RECT 139.525 207.000 140.735 207.750 ;
        RECT 141.540 207.720 141.710 207.910 ;
        RECT 141.965 207.745 142.135 208.475 ;
        RECT 142.310 208.400 142.570 209.550 ;
        RECT 142.835 208.620 143.005 209.380 ;
        RECT 143.220 208.790 143.550 209.550 ;
        RECT 142.835 208.450 143.550 208.620 ;
        RECT 143.720 208.475 143.975 209.380 ;
        RECT 142.745 207.900 143.100 208.270 ;
        RECT 143.380 208.240 143.550 208.450 ;
        RECT 143.380 207.910 143.635 208.240 ;
        RECT 140.995 207.550 141.710 207.720 ;
        RECT 140.995 207.170 141.165 207.550 ;
        RECT 141.380 207.000 141.710 207.380 ;
        RECT 141.880 207.170 142.135 207.745 ;
        RECT 142.310 207.000 142.570 207.840 ;
        RECT 143.380 207.720 143.550 207.910 ;
        RECT 143.805 207.745 143.975 208.475 ;
        RECT 144.150 208.400 144.410 209.550 ;
        RECT 144.675 208.620 144.845 209.380 ;
        RECT 145.060 208.790 145.390 209.550 ;
        RECT 144.675 208.450 145.390 208.620 ;
        RECT 145.560 208.475 145.815 209.380 ;
        RECT 144.585 207.900 144.940 208.270 ;
        RECT 145.220 208.240 145.390 208.450 ;
        RECT 145.220 207.910 145.475 208.240 ;
        RECT 142.835 207.550 143.550 207.720 ;
        RECT 142.835 207.170 143.005 207.550 ;
        RECT 143.220 207.000 143.550 207.380 ;
        RECT 143.720 207.170 143.975 207.745 ;
        RECT 144.150 207.000 144.410 207.840 ;
        RECT 145.220 207.720 145.390 207.910 ;
        RECT 145.645 207.745 145.815 208.475 ;
        RECT 145.990 208.400 146.250 209.550 ;
        RECT 146.425 208.460 147.635 209.550 ;
        RECT 146.425 207.920 146.945 208.460 ;
        RECT 144.675 207.550 145.390 207.720 ;
        RECT 144.675 207.170 144.845 207.550 ;
        RECT 145.060 207.000 145.390 207.380 ;
        RECT 145.560 207.170 145.815 207.745 ;
        RECT 145.990 207.000 146.250 207.840 ;
        RECT 147.115 207.750 147.635 208.290 ;
        RECT 146.425 207.000 147.635 207.750 ;
        RECT 13.860 206.830 147.720 207.000 ;
        RECT 13.945 206.080 15.155 206.830 ;
        RECT 13.945 205.540 14.465 206.080 ;
        RECT 15.330 205.990 15.590 206.830 ;
        RECT 15.765 206.085 16.020 206.660 ;
        RECT 16.190 206.450 16.520 206.830 ;
        RECT 16.735 206.280 16.905 206.660 ;
        RECT 16.190 206.110 16.905 206.280 ;
        RECT 14.635 205.370 15.155 205.910 ;
        RECT 13.945 204.280 15.155 205.370 ;
        RECT 15.330 204.280 15.590 205.430 ;
        RECT 15.765 205.355 15.935 206.085 ;
        RECT 16.190 205.920 16.360 206.110 ;
        RECT 17.170 205.990 17.430 206.830 ;
        RECT 17.605 206.085 17.860 206.660 ;
        RECT 18.030 206.450 18.360 206.830 ;
        RECT 18.575 206.280 18.745 206.660 ;
        RECT 18.030 206.110 18.745 206.280 ;
        RECT 19.005 206.155 19.265 206.660 ;
        RECT 19.445 206.450 19.775 206.830 ;
        RECT 19.955 206.280 20.125 206.660 ;
        RECT 16.105 205.590 16.360 205.920 ;
        RECT 16.190 205.380 16.360 205.590 ;
        RECT 16.640 205.560 16.995 205.930 ;
        RECT 15.765 204.450 16.020 205.355 ;
        RECT 16.190 205.210 16.905 205.380 ;
        RECT 16.190 204.280 16.520 205.040 ;
        RECT 16.735 204.450 16.905 205.210 ;
        RECT 17.170 204.280 17.430 205.430 ;
        RECT 17.605 205.355 17.775 206.085 ;
        RECT 18.030 205.920 18.200 206.110 ;
        RECT 17.945 205.590 18.200 205.920 ;
        RECT 18.030 205.380 18.200 205.590 ;
        RECT 18.480 205.560 18.835 205.930 ;
        RECT 17.605 204.450 17.860 205.355 ;
        RECT 18.030 205.210 18.745 205.380 ;
        RECT 18.030 204.280 18.360 205.040 ;
        RECT 18.575 204.450 18.745 205.210 ;
        RECT 19.005 205.355 19.175 206.155 ;
        RECT 19.460 206.110 20.125 206.280 ;
        RECT 19.460 205.855 19.630 206.110 ;
        RECT 20.385 206.060 23.895 206.830 ;
        RECT 19.345 205.525 19.630 205.855 ;
        RECT 19.865 205.560 20.195 205.930 ;
        RECT 20.385 205.540 22.035 206.060 ;
        RECT 24.535 206.020 24.805 206.830 ;
        RECT 24.975 206.020 25.305 206.660 ;
        RECT 25.475 206.020 25.715 206.830 ;
        RECT 26.105 206.200 26.435 206.560 ;
        RECT 27.055 206.370 27.305 206.830 ;
        RECT 27.475 206.370 28.035 206.660 ;
        RECT 19.460 205.380 19.630 205.525 ;
        RECT 19.005 204.450 19.275 205.355 ;
        RECT 19.460 205.210 20.125 205.380 ;
        RECT 22.205 205.370 23.895 205.890 ;
        RECT 24.525 205.590 24.875 205.840 ;
        RECT 25.045 205.420 25.215 206.020 ;
        RECT 26.105 206.010 27.495 206.200 ;
        RECT 27.325 205.920 27.495 206.010 ;
        RECT 25.385 205.590 25.735 205.840 ;
        RECT 25.920 205.590 26.595 205.840 ;
        RECT 26.815 205.590 27.155 205.840 ;
        RECT 27.325 205.590 27.615 205.920 ;
        RECT 19.445 204.280 19.775 205.040 ;
        RECT 19.955 204.450 20.125 205.210 ;
        RECT 20.385 204.280 23.895 205.370 ;
        RECT 24.535 204.280 24.865 205.420 ;
        RECT 25.045 205.250 25.725 205.420 ;
        RECT 25.395 204.465 25.725 205.250 ;
        RECT 25.920 205.230 26.185 205.590 ;
        RECT 27.325 205.340 27.495 205.590 ;
        RECT 26.555 205.170 27.495 205.340 ;
        RECT 26.105 204.280 26.385 204.950 ;
        RECT 26.555 204.620 26.855 205.170 ;
        RECT 27.785 205.000 28.035 206.370 ;
        RECT 28.665 206.010 28.925 206.830 ;
        RECT 29.095 206.010 29.425 206.430 ;
        RECT 29.605 206.260 29.865 206.660 ;
        RECT 30.035 206.430 30.365 206.830 ;
        RECT 30.535 206.260 30.705 206.610 ;
        RECT 30.875 206.430 31.250 206.830 ;
        RECT 29.605 206.090 31.270 206.260 ;
        RECT 31.440 206.155 31.715 206.500 ;
        RECT 29.175 205.920 29.425 206.010 ;
        RECT 31.100 205.920 31.270 206.090 ;
        RECT 28.670 205.590 29.005 205.840 ;
        RECT 29.175 205.590 29.890 205.920 ;
        RECT 30.105 205.590 30.930 205.920 ;
        RECT 31.100 205.590 31.375 205.920 ;
        RECT 27.055 204.280 27.385 205.000 ;
        RECT 27.575 204.450 28.035 205.000 ;
        RECT 28.665 204.280 28.925 205.420 ;
        RECT 29.175 205.030 29.345 205.590 ;
        RECT 29.605 205.130 29.935 205.420 ;
        RECT 30.105 205.300 30.350 205.590 ;
        RECT 31.100 205.420 31.270 205.590 ;
        RECT 31.545 205.420 31.715 206.155 ;
        RECT 31.885 206.030 32.580 206.660 ;
        RECT 32.785 206.030 33.095 206.830 ;
        RECT 33.265 206.060 34.935 206.830 ;
        RECT 31.905 205.590 32.240 205.840 ;
        RECT 32.410 205.430 32.580 206.030 ;
        RECT 32.750 205.590 33.085 205.860 ;
        RECT 33.265 205.540 34.015 206.060 ;
        RECT 35.105 206.030 35.800 206.660 ;
        RECT 36.005 206.030 36.315 206.830 ;
        RECT 30.610 205.250 31.270 205.420 ;
        RECT 30.610 205.130 30.780 205.250 ;
        RECT 29.605 204.960 30.780 205.130 ;
        RECT 29.165 204.460 30.780 204.790 ;
        RECT 30.950 204.280 31.230 205.080 ;
        RECT 31.440 204.450 31.715 205.420 ;
        RECT 31.885 204.280 32.145 205.420 ;
        RECT 32.315 204.450 32.645 205.430 ;
        RECT 32.815 204.280 33.095 205.420 ;
        RECT 34.185 205.370 34.935 205.890 ;
        RECT 35.125 205.590 35.460 205.840 ;
        RECT 35.630 205.430 35.800 206.030 ;
        RECT 36.525 206.010 36.755 206.830 ;
        RECT 36.925 206.030 37.255 206.660 ;
        RECT 35.970 205.590 36.305 205.860 ;
        RECT 36.505 205.590 36.835 205.840 ;
        RECT 37.005 205.430 37.255 206.030 ;
        RECT 37.425 206.010 37.635 206.830 ;
        RECT 37.870 206.430 38.205 206.830 ;
        RECT 38.375 206.260 38.580 206.660 ;
        RECT 38.790 206.350 39.065 206.830 ;
        RECT 39.275 206.330 39.535 206.660 ;
        RECT 37.895 206.090 38.580 206.260 ;
        RECT 33.265 204.280 34.935 205.370 ;
        RECT 35.105 204.280 35.365 205.420 ;
        RECT 35.535 204.450 35.865 205.430 ;
        RECT 36.035 204.280 36.315 205.420 ;
        RECT 36.525 204.280 36.755 205.420 ;
        RECT 36.925 204.450 37.255 205.430 ;
        RECT 37.425 204.280 37.635 205.420 ;
        RECT 37.895 205.060 38.235 206.090 ;
        RECT 38.405 205.420 38.655 205.920 ;
        RECT 38.835 205.590 39.195 206.170 ;
        RECT 39.365 205.420 39.535 206.330 ;
        RECT 39.705 206.105 39.995 206.830 ;
        RECT 40.165 206.070 40.875 206.660 ;
        RECT 41.385 206.300 41.715 206.660 ;
        RECT 41.915 206.470 42.245 206.830 ;
        RECT 42.415 206.300 42.745 206.660 ;
        RECT 41.385 206.090 42.745 206.300 ;
        RECT 42.935 206.105 43.265 206.615 ;
        RECT 43.435 206.430 43.765 206.830 ;
        RECT 44.815 206.260 45.145 206.600 ;
        RECT 45.315 206.430 45.645 206.830 ;
        RECT 46.605 206.430 47.195 206.660 ;
        RECT 48.240 206.430 48.570 206.830 ;
        RECT 38.405 205.250 39.535 205.420 ;
        RECT 37.895 204.885 38.560 205.060 ;
        RECT 37.870 204.280 38.205 204.705 ;
        RECT 38.375 204.480 38.560 204.885 ;
        RECT 38.765 204.280 39.095 205.060 ;
        RECT 39.265 204.480 39.535 205.250 ;
        RECT 39.705 204.280 39.995 205.445 ;
        RECT 40.165 205.130 40.370 206.070 ;
        RECT 40.540 205.300 40.870 205.840 ;
        RECT 41.045 205.590 41.540 205.920 ;
        RECT 41.860 205.590 42.235 205.920 ;
        RECT 42.445 205.590 42.755 205.920 ;
        RECT 41.045 205.300 41.370 205.590 ;
        RECT 40.165 205.100 40.395 205.130 ;
        RECT 41.565 205.100 41.895 205.320 ;
        RECT 40.165 204.870 41.895 205.100 ;
        RECT 40.165 204.450 40.865 204.870 ;
        RECT 41.065 204.280 41.395 204.640 ;
        RECT 41.565 204.470 41.895 204.870 ;
        RECT 42.065 204.620 42.235 205.590 ;
        RECT 42.935 205.470 43.125 206.105 ;
        RECT 43.435 206.090 45.800 206.260 ;
        RECT 43.435 205.920 43.605 206.090 ;
        RECT 43.295 205.590 43.605 205.920 ;
        RECT 43.775 205.590 44.080 205.920 ;
        RECT 42.935 205.340 43.155 205.470 ;
        RECT 42.415 204.280 42.745 205.340 ;
        RECT 42.935 204.490 43.265 205.340 ;
        RECT 43.435 204.280 43.685 205.420 ;
        RECT 43.865 205.260 44.080 205.590 ;
        RECT 44.255 205.260 44.540 205.920 ;
        RECT 44.735 205.260 45.000 205.920 ;
        RECT 45.215 205.260 45.460 205.920 ;
        RECT 45.630 205.090 45.800 206.090 ;
        RECT 43.875 204.920 45.165 205.090 ;
        RECT 43.875 204.500 44.125 204.920 ;
        RECT 44.355 204.280 44.685 204.750 ;
        RECT 44.915 204.500 45.165 204.920 ;
        RECT 45.345 204.920 45.800 205.090 ;
        RECT 46.605 205.420 46.895 206.430 ;
        RECT 48.770 206.260 49.195 206.470 ;
        RECT 47.065 206.090 49.195 206.260 ;
        RECT 47.065 205.590 47.235 206.090 ;
        RECT 47.525 205.590 47.855 205.920 ;
        RECT 48.045 205.590 48.315 205.920 ;
        RECT 48.505 205.590 48.855 205.920 ;
        RECT 46.605 205.250 48.150 205.420 ;
        RECT 45.345 204.490 45.675 204.920 ;
        RECT 46.605 204.450 47.195 205.250 ;
        RECT 47.365 204.280 47.650 205.080 ;
        RECT 47.820 204.450 48.150 205.250 ;
        RECT 48.320 204.280 48.570 205.420 ;
        RECT 49.025 205.320 49.195 206.090 ;
        RECT 50.285 206.030 50.595 206.830 ;
        RECT 50.800 206.030 51.495 206.660 ;
        RECT 52.170 206.370 52.920 206.660 ;
        RECT 53.430 206.370 53.760 206.830 ;
        RECT 50.295 205.590 50.630 205.860 ;
        RECT 50.800 205.430 50.970 206.030 ;
        RECT 51.140 205.590 51.475 205.840 ;
        RECT 48.770 204.990 49.195 205.320 ;
        RECT 50.285 204.280 50.565 205.420 ;
        RECT 50.735 204.450 51.065 205.430 ;
        RECT 51.235 204.280 51.495 205.420 ;
        RECT 52.170 205.080 52.540 206.370 ;
        RECT 53.980 206.180 54.250 206.390 ;
        RECT 52.915 206.010 54.250 206.180 ;
        RECT 54.515 206.180 54.685 206.660 ;
        RECT 54.855 206.350 55.185 206.830 ;
        RECT 55.410 206.410 56.945 206.660 ;
        RECT 55.410 206.180 55.580 206.410 ;
        RECT 54.515 206.010 55.580 206.180 ;
        RECT 52.915 205.840 53.085 206.010 ;
        RECT 55.760 205.840 56.040 206.240 ;
        RECT 52.710 205.590 53.085 205.840 ;
        RECT 53.255 205.600 53.730 205.840 ;
        RECT 53.900 205.600 54.250 205.840 ;
        RECT 54.430 205.630 54.780 205.840 ;
        RECT 54.950 205.640 55.395 205.840 ;
        RECT 55.565 205.640 56.040 205.840 ;
        RECT 56.310 205.840 56.595 206.240 ;
        RECT 56.775 206.180 56.945 206.410 ;
        RECT 57.115 206.350 57.445 206.830 ;
        RECT 57.660 206.330 57.915 206.660 ;
        RECT 57.705 206.320 57.915 206.330 ;
        RECT 57.730 206.250 57.915 206.320 ;
        RECT 56.775 206.010 57.575 206.180 ;
        RECT 56.310 205.640 56.640 205.840 ;
        RECT 56.810 205.640 57.175 205.840 ;
        RECT 52.915 205.420 53.085 205.590 ;
        RECT 57.405 205.460 57.575 206.010 ;
        RECT 52.915 205.250 54.250 205.420 ;
        RECT 53.970 205.090 54.250 205.250 ;
        RECT 54.515 205.290 57.575 205.460 ;
        RECT 52.170 204.910 53.340 205.080 ;
        RECT 52.625 204.280 52.840 204.740 ;
        RECT 53.010 204.450 53.340 204.910 ;
        RECT 53.510 204.280 53.760 205.080 ;
        RECT 54.515 204.450 54.685 205.290 ;
        RECT 57.745 205.120 57.915 206.250 ;
        RECT 54.855 204.620 55.185 205.120 ;
        RECT 55.355 204.880 56.990 205.120 ;
        RECT 55.355 204.790 55.585 204.880 ;
        RECT 55.695 204.620 56.025 204.660 ;
        RECT 54.855 204.450 56.025 204.620 ;
        RECT 56.215 204.280 56.570 204.700 ;
        RECT 56.740 204.450 56.990 204.880 ;
        RECT 57.160 204.280 57.490 205.040 ;
        RECT 57.660 204.450 57.915 205.120 ;
        RECT 58.105 206.330 58.365 206.660 ;
        RECT 58.535 206.470 58.865 206.830 ;
        RECT 59.120 206.450 60.420 206.660 ;
        RECT 58.105 206.320 58.335 206.330 ;
        RECT 58.105 205.130 58.275 206.320 ;
        RECT 59.120 206.300 59.290 206.450 ;
        RECT 58.535 206.175 59.290 206.300 ;
        RECT 58.445 206.130 59.290 206.175 ;
        RECT 58.445 206.010 58.715 206.130 ;
        RECT 58.445 205.435 58.615 206.010 ;
        RECT 58.845 205.570 59.255 205.875 ;
        RECT 59.545 205.840 59.755 206.240 ;
        RECT 59.425 205.630 59.755 205.840 ;
        RECT 60.000 205.840 60.220 206.240 ;
        RECT 60.695 206.065 61.150 206.830 ;
        RECT 61.985 206.200 62.315 206.560 ;
        RECT 62.935 206.370 63.185 206.830 ;
        RECT 63.355 206.370 63.915 206.660 ;
        RECT 61.985 206.010 63.375 206.200 ;
        RECT 63.205 205.920 63.375 206.010 ;
        RECT 60.000 205.630 60.475 205.840 ;
        RECT 60.665 205.640 61.155 205.840 ;
        RECT 61.800 205.590 62.475 205.840 ;
        RECT 62.695 205.590 63.035 205.840 ;
        RECT 63.205 205.590 63.495 205.920 ;
        RECT 58.445 205.400 58.645 205.435 ;
        RECT 59.975 205.400 61.150 205.460 ;
        RECT 58.445 205.290 61.150 205.400 ;
        RECT 58.505 205.230 60.305 205.290 ;
        RECT 59.975 205.200 60.305 205.230 ;
        RECT 58.105 204.450 58.365 205.130 ;
        RECT 58.535 204.280 58.785 205.060 ;
        RECT 59.035 205.030 59.870 205.040 ;
        RECT 60.460 205.030 60.645 205.120 ;
        RECT 59.035 204.830 60.645 205.030 ;
        RECT 59.035 204.450 59.285 204.830 ;
        RECT 60.415 204.790 60.645 204.830 ;
        RECT 60.895 204.670 61.150 205.290 ;
        RECT 61.800 205.230 62.065 205.590 ;
        RECT 63.205 205.340 63.375 205.590 ;
        RECT 62.435 205.170 63.375 205.340 ;
        RECT 59.455 204.280 59.810 204.660 ;
        RECT 60.815 204.450 61.150 204.670 ;
        RECT 61.985 204.280 62.265 204.950 ;
        RECT 62.435 204.620 62.735 205.170 ;
        RECT 63.665 205.000 63.915 206.370 ;
        RECT 64.085 206.030 64.395 206.830 ;
        RECT 64.600 206.030 65.295 206.660 ;
        RECT 65.465 206.105 65.755 206.830 ;
        RECT 65.930 206.090 66.185 206.660 ;
        RECT 66.355 206.430 66.685 206.830 ;
        RECT 67.110 206.295 67.640 206.660 ;
        RECT 67.110 206.260 67.285 206.295 ;
        RECT 66.355 206.090 67.285 206.260 ;
        RECT 67.830 206.150 68.105 206.660 ;
        RECT 64.600 205.980 64.775 206.030 ;
        RECT 64.095 205.590 64.430 205.860 ;
        RECT 64.600 205.430 64.770 205.980 ;
        RECT 64.940 205.590 65.275 205.840 ;
        RECT 62.935 204.280 63.265 205.000 ;
        RECT 63.455 204.450 63.915 205.000 ;
        RECT 64.085 204.280 64.365 205.420 ;
        RECT 64.535 204.450 64.865 205.430 ;
        RECT 65.035 204.280 65.295 205.420 ;
        RECT 65.465 204.280 65.755 205.445 ;
        RECT 65.930 205.420 66.100 206.090 ;
        RECT 66.355 205.920 66.525 206.090 ;
        RECT 66.270 205.590 66.525 205.920 ;
        RECT 66.750 205.590 66.945 205.920 ;
        RECT 65.930 204.450 66.265 205.420 ;
        RECT 66.435 204.280 66.605 205.420 ;
        RECT 66.775 204.620 66.945 205.590 ;
        RECT 67.115 204.960 67.285 206.090 ;
        RECT 67.455 205.300 67.625 206.100 ;
        RECT 67.825 205.980 68.105 206.150 ;
        RECT 67.830 205.500 68.105 205.980 ;
        RECT 68.275 205.300 68.465 206.660 ;
        RECT 68.645 206.295 69.155 206.830 ;
        RECT 69.375 206.020 69.620 206.625 ;
        RECT 70.065 206.030 70.760 206.660 ;
        RECT 70.965 206.030 71.275 206.830 ;
        RECT 71.445 206.070 72.155 206.660 ;
        RECT 72.665 206.300 72.995 206.660 ;
        RECT 73.195 206.470 73.525 206.830 ;
        RECT 73.695 206.300 74.025 206.660 ;
        RECT 74.295 206.350 74.595 206.830 ;
        RECT 72.665 206.090 74.025 206.300 ;
        RECT 74.765 206.180 75.025 206.635 ;
        RECT 75.195 206.350 75.455 206.830 ;
        RECT 75.635 206.180 75.895 206.635 ;
        RECT 76.065 206.350 76.315 206.830 ;
        RECT 76.495 206.180 76.755 206.635 ;
        RECT 76.925 206.350 77.175 206.830 ;
        RECT 77.355 206.180 77.615 206.635 ;
        RECT 77.785 206.350 78.030 206.830 ;
        RECT 78.200 206.180 78.475 206.635 ;
        RECT 78.645 206.350 78.890 206.830 ;
        RECT 79.060 206.180 79.320 206.635 ;
        RECT 79.490 206.350 79.750 206.830 ;
        RECT 79.920 206.180 80.180 206.635 ;
        RECT 80.350 206.350 80.610 206.830 ;
        RECT 80.780 206.180 81.040 206.635 ;
        RECT 81.210 206.270 81.470 206.830 ;
        RECT 68.665 205.850 69.895 206.020 ;
        RECT 70.585 205.980 70.760 206.030 ;
        RECT 67.455 205.130 68.465 205.300 ;
        RECT 68.635 205.285 69.385 205.475 ;
        RECT 67.115 204.790 68.240 204.960 ;
        RECT 68.635 204.620 68.805 205.285 ;
        RECT 69.555 205.040 69.895 205.850 ;
        RECT 70.085 205.590 70.420 205.840 ;
        RECT 70.590 205.430 70.760 205.980 ;
        RECT 71.445 205.980 71.675 206.070 ;
        RECT 74.295 206.010 81.040 206.180 ;
        RECT 70.930 205.590 71.265 205.860 ;
        RECT 66.775 204.450 68.805 204.620 ;
        RECT 68.975 204.280 69.145 205.040 ;
        RECT 69.380 204.630 69.895 205.040 ;
        RECT 70.065 204.280 70.325 205.420 ;
        RECT 70.495 204.450 70.825 205.430 ;
        RECT 70.995 204.280 71.275 205.420 ;
        RECT 71.445 205.100 71.650 205.980 ;
        RECT 71.820 205.300 72.150 205.840 ;
        RECT 72.325 205.590 72.820 205.920 ;
        RECT 73.140 205.590 73.515 205.920 ;
        RECT 73.725 205.590 74.035 205.920 ;
        RECT 72.325 205.300 72.650 205.590 ;
        RECT 72.845 205.100 73.175 205.320 ;
        RECT 71.445 204.870 73.175 205.100 ;
        RECT 71.445 204.450 72.145 204.870 ;
        RECT 72.345 204.280 72.675 204.640 ;
        RECT 72.845 204.470 73.175 204.870 ;
        RECT 73.345 204.620 73.515 205.590 ;
        RECT 74.295 205.420 75.460 206.010 ;
        RECT 81.640 205.840 81.890 206.650 ;
        RECT 82.070 206.305 82.330 206.830 ;
        RECT 82.500 205.840 82.750 206.650 ;
        RECT 82.930 206.320 83.235 206.830 ;
        RECT 75.630 205.590 82.750 205.840 ;
        RECT 82.920 205.590 83.235 206.150 ;
        RECT 83.425 206.140 83.665 206.660 ;
        RECT 83.835 206.335 84.230 206.830 ;
        RECT 84.795 206.500 84.965 206.645 ;
        RECT 84.590 206.305 84.965 206.500 ;
        RECT 73.695 204.280 74.025 205.340 ;
        RECT 74.295 205.195 81.040 205.420 ;
        RECT 74.295 204.280 74.565 205.025 ;
        RECT 74.735 204.455 75.025 205.195 ;
        RECT 75.635 205.180 81.040 205.195 ;
        RECT 75.195 204.285 75.450 205.010 ;
        RECT 75.635 204.455 75.895 205.180 ;
        RECT 76.065 204.285 76.310 205.010 ;
        RECT 76.495 204.455 76.755 205.180 ;
        RECT 76.925 204.285 77.170 205.010 ;
        RECT 77.355 204.455 77.615 205.180 ;
        RECT 77.785 204.285 78.030 205.010 ;
        RECT 78.200 204.455 78.460 205.180 ;
        RECT 78.630 204.285 78.890 205.010 ;
        RECT 79.060 204.455 79.320 205.180 ;
        RECT 79.490 204.285 79.750 205.010 ;
        RECT 79.920 204.455 80.180 205.180 ;
        RECT 80.350 204.285 80.610 205.010 ;
        RECT 80.780 204.455 81.040 205.180 ;
        RECT 81.210 204.285 81.470 205.080 ;
        RECT 81.640 204.455 81.890 205.590 ;
        RECT 75.195 204.280 81.470 204.285 ;
        RECT 82.070 204.280 82.330 205.090 ;
        RECT 82.505 204.450 82.750 205.590 ;
        RECT 83.425 205.470 83.600 206.140 ;
        RECT 84.590 205.970 84.760 206.305 ;
        RECT 85.245 206.260 85.485 206.635 ;
        RECT 85.655 206.325 85.990 206.830 ;
        RECT 85.245 206.110 85.465 206.260 ;
        RECT 83.775 205.610 84.760 205.970 ;
        RECT 84.930 205.780 85.465 206.110 ;
        RECT 83.775 205.590 85.060 205.610 ;
        RECT 83.425 205.335 83.635 205.470 ;
        RECT 84.200 205.440 85.060 205.590 ;
        RECT 82.930 204.280 83.225 205.090 ;
        RECT 83.425 204.550 83.730 205.335 ;
        RECT 83.905 204.960 84.600 205.270 ;
        RECT 83.910 204.280 84.595 204.750 ;
        RECT 84.775 204.495 85.060 205.440 ;
        RECT 85.230 205.130 85.465 205.780 ;
        RECT 85.635 205.300 85.935 206.150 ;
        RECT 86.165 206.030 86.475 206.830 ;
        RECT 86.680 206.030 87.375 206.660 ;
        RECT 88.485 206.140 88.725 206.660 ;
        RECT 88.895 206.335 89.290 206.830 ;
        RECT 89.855 206.500 90.025 206.645 ;
        RECT 89.650 206.305 90.025 206.500 ;
        RECT 86.175 205.590 86.510 205.860 ;
        RECT 86.680 205.430 86.850 206.030 ;
        RECT 87.020 205.590 87.355 205.840 ;
        RECT 88.485 205.470 88.660 206.140 ;
        RECT 89.650 205.970 89.820 206.305 ;
        RECT 90.305 206.260 90.545 206.635 ;
        RECT 90.715 206.325 91.050 206.830 ;
        RECT 90.305 206.110 90.525 206.260 ;
        RECT 88.835 205.610 89.820 205.970 ;
        RECT 89.990 205.780 90.525 206.110 ;
        RECT 88.835 205.590 90.120 205.610 ;
        RECT 85.230 204.900 85.905 205.130 ;
        RECT 85.235 204.280 85.565 204.730 ;
        RECT 85.735 204.470 85.905 204.900 ;
        RECT 86.165 204.280 86.445 205.420 ;
        RECT 86.615 204.450 86.945 205.430 ;
        RECT 87.115 204.280 87.375 205.420 ;
        RECT 88.485 205.335 88.695 205.470 ;
        RECT 89.260 205.440 90.120 205.590 ;
        RECT 88.485 204.550 88.790 205.335 ;
        RECT 88.965 204.960 89.660 205.270 ;
        RECT 88.970 204.280 89.655 204.750 ;
        RECT 89.835 204.495 90.120 205.440 ;
        RECT 90.290 205.130 90.525 205.780 ;
        RECT 90.695 205.300 90.995 206.150 ;
        RECT 91.225 206.105 91.515 206.830 ;
        RECT 91.745 206.010 91.955 206.830 ;
        RECT 92.125 206.030 92.455 206.660 ;
        RECT 90.290 204.900 90.965 205.130 ;
        RECT 90.295 204.280 90.625 204.730 ;
        RECT 90.795 204.470 90.965 204.900 ;
        RECT 91.225 204.280 91.515 205.445 ;
        RECT 92.125 205.430 92.375 206.030 ;
        RECT 92.625 206.010 92.855 206.830 ;
        RECT 93.065 206.060 94.735 206.830 ;
        RECT 92.545 205.590 92.875 205.840 ;
        RECT 93.065 205.540 93.815 206.060 ;
        RECT 94.905 206.030 95.600 206.660 ;
        RECT 95.805 206.030 96.115 206.830 ;
        RECT 96.290 206.090 96.545 206.660 ;
        RECT 96.715 206.430 97.045 206.830 ;
        RECT 97.470 206.295 98.000 206.660 ;
        RECT 97.470 206.260 97.645 206.295 ;
        RECT 96.715 206.090 97.645 206.260 ;
        RECT 91.745 204.280 91.955 205.420 ;
        RECT 92.125 204.450 92.455 205.430 ;
        RECT 92.625 204.280 92.855 205.420 ;
        RECT 93.985 205.370 94.735 205.890 ;
        RECT 94.925 205.590 95.260 205.840 ;
        RECT 95.430 205.430 95.600 206.030 ;
        RECT 95.770 205.590 96.105 205.860 ;
        RECT 93.065 204.280 94.735 205.370 ;
        RECT 94.905 204.280 95.165 205.420 ;
        RECT 95.335 204.450 95.665 205.430 ;
        RECT 96.290 205.420 96.460 206.090 ;
        RECT 96.715 205.920 96.885 206.090 ;
        RECT 96.630 205.590 96.885 205.920 ;
        RECT 97.110 205.590 97.305 205.920 ;
        RECT 95.835 204.280 96.115 205.420 ;
        RECT 96.290 204.450 96.625 205.420 ;
        RECT 96.795 204.280 96.965 205.420 ;
        RECT 97.135 204.620 97.305 205.590 ;
        RECT 97.475 204.960 97.645 206.090 ;
        RECT 97.815 205.300 97.985 206.100 ;
        RECT 98.190 205.810 98.465 206.660 ;
        RECT 98.185 205.640 98.465 205.810 ;
        RECT 98.190 205.500 98.465 205.640 ;
        RECT 98.635 205.300 98.825 206.660 ;
        RECT 99.005 206.295 99.515 206.830 ;
        RECT 99.735 206.020 99.980 206.625 ;
        RECT 100.435 206.105 100.765 206.615 ;
        RECT 100.935 206.430 101.265 206.830 ;
        RECT 102.315 206.260 102.645 206.600 ;
        RECT 102.815 206.430 103.145 206.830 ;
        RECT 103.645 206.260 104.070 206.470 ;
        RECT 104.270 206.430 104.600 206.830 ;
        RECT 105.645 206.430 106.235 206.660 ;
        RECT 99.025 205.850 100.255 206.020 ;
        RECT 97.815 205.130 98.825 205.300 ;
        RECT 98.995 205.285 99.745 205.475 ;
        RECT 97.475 204.790 98.600 204.960 ;
        RECT 98.995 204.620 99.165 205.285 ;
        RECT 99.915 205.040 100.255 205.850 ;
        RECT 97.135 204.450 99.165 204.620 ;
        RECT 99.335 204.280 99.505 205.040 ;
        RECT 99.740 204.630 100.255 205.040 ;
        RECT 100.435 205.340 100.625 206.105 ;
        RECT 100.935 206.090 103.300 206.260 ;
        RECT 100.935 205.920 101.105 206.090 ;
        RECT 100.795 205.590 101.105 205.920 ;
        RECT 101.275 205.590 101.580 205.920 ;
        RECT 100.435 204.490 100.765 205.340 ;
        RECT 100.935 204.280 101.185 205.420 ;
        RECT 101.365 205.260 101.580 205.590 ;
        RECT 101.755 205.260 102.040 205.920 ;
        RECT 102.235 205.260 102.500 205.920 ;
        RECT 102.715 205.260 102.960 205.920 ;
        RECT 103.130 205.090 103.300 206.090 ;
        RECT 101.375 204.920 102.665 205.090 ;
        RECT 101.375 204.500 101.625 204.920 ;
        RECT 101.855 204.280 102.185 204.750 ;
        RECT 102.415 204.500 102.665 204.920 ;
        RECT 102.845 204.920 103.300 205.090 ;
        RECT 103.645 206.090 105.775 206.260 ;
        RECT 103.645 205.320 103.815 206.090 ;
        RECT 103.985 205.590 104.335 205.920 ;
        RECT 104.525 205.590 104.795 205.920 ;
        RECT 104.985 205.590 105.315 205.920 ;
        RECT 105.605 205.590 105.775 206.090 ;
        RECT 105.945 205.420 106.235 206.430 ;
        RECT 106.870 206.325 107.205 206.830 ;
        RECT 107.375 206.260 107.615 206.635 ;
        RECT 107.895 206.500 108.065 206.645 ;
        RECT 107.895 206.305 108.270 206.500 ;
        RECT 108.630 206.335 109.025 206.830 ;
        RECT 103.645 204.990 104.070 205.320 ;
        RECT 102.845 204.490 103.175 204.920 ;
        RECT 104.270 204.280 104.520 205.420 ;
        RECT 104.690 205.250 106.235 205.420 ;
        RECT 106.925 205.300 107.225 206.150 ;
        RECT 107.395 206.110 107.615 206.260 ;
        RECT 107.395 205.780 107.930 206.110 ;
        RECT 108.100 205.970 108.270 206.305 ;
        RECT 109.195 206.140 109.435 206.660 ;
        RECT 104.690 204.450 105.020 205.250 ;
        RECT 105.190 204.280 105.475 205.080 ;
        RECT 105.645 204.450 106.235 205.250 ;
        RECT 107.395 205.130 107.630 205.780 ;
        RECT 108.100 205.610 109.085 205.970 ;
        RECT 106.955 204.900 107.630 205.130 ;
        RECT 107.800 205.590 109.085 205.610 ;
        RECT 107.800 205.440 108.660 205.590 ;
        RECT 106.955 204.470 107.125 204.900 ;
        RECT 107.295 204.280 107.625 204.730 ;
        RECT 107.800 204.495 108.085 205.440 ;
        RECT 109.260 205.335 109.435 206.140 ;
        RECT 108.260 204.960 108.955 205.270 ;
        RECT 108.265 204.280 108.950 204.750 ;
        RECT 109.130 204.550 109.435 205.335 ;
        RECT 109.625 206.355 109.965 206.615 ;
        RECT 109.625 204.750 109.885 206.355 ;
        RECT 110.135 206.350 110.465 206.830 ;
        RECT 110.655 206.180 111.070 206.615 ;
        RECT 111.240 206.315 112.190 206.500 ;
        RECT 110.055 206.105 111.070 206.180 ;
        RECT 110.055 206.010 110.875 206.105 ;
        RECT 110.055 205.090 110.225 206.010 ;
        RECT 110.545 205.280 110.875 205.840 ;
        RECT 111.075 205.590 111.455 205.920 ;
        RECT 111.765 205.590 111.985 206.315 ;
        RECT 112.420 205.920 112.625 206.520 ;
        RECT 112.795 206.105 113.135 206.830 ;
        RECT 113.305 206.155 113.580 206.500 ;
        RECT 113.770 206.430 114.145 206.830 ;
        RECT 114.315 206.260 114.485 206.610 ;
        RECT 114.655 206.430 114.985 206.830 ;
        RECT 115.155 206.260 115.415 206.660 ;
        RECT 111.075 205.470 111.375 205.590 ;
        RECT 111.065 205.300 111.375 205.470 ;
        RECT 111.075 205.295 111.375 205.300 ;
        RECT 112.245 205.290 112.625 205.920 ;
        RECT 112.855 205.290 113.110 205.920 ;
        RECT 113.305 205.420 113.475 206.155 ;
        RECT 113.750 206.090 115.415 206.260 ;
        RECT 113.750 205.920 113.920 206.090 ;
        RECT 115.595 206.010 115.925 206.430 ;
        RECT 116.095 206.010 116.355 206.830 ;
        RECT 116.985 206.105 117.275 206.830 ;
        RECT 117.445 206.330 117.785 206.830 ;
        RECT 115.595 205.920 115.845 206.010 ;
        RECT 113.645 205.590 113.920 205.920 ;
        RECT 114.090 205.590 114.915 205.920 ;
        RECT 115.130 205.590 115.845 205.920 ;
        RECT 116.015 205.590 116.350 205.840 ;
        RECT 117.445 205.590 117.785 206.160 ;
        RECT 117.955 205.920 118.200 206.610 ;
        RECT 118.395 206.330 118.725 206.830 ;
        RECT 118.925 206.260 119.095 206.610 ;
        RECT 119.270 206.430 119.600 206.830 ;
        RECT 119.770 206.260 119.940 206.610 ;
        RECT 120.110 206.430 120.490 206.830 ;
        RECT 118.925 206.090 120.510 206.260 ;
        RECT 120.680 206.155 120.955 206.500 ;
        RECT 120.340 205.920 120.510 206.090 ;
        RECT 117.955 205.590 118.610 205.920 ;
        RECT 113.750 205.420 113.920 205.590 ;
        RECT 110.055 204.920 110.905 205.090 ;
        RECT 109.625 204.490 109.965 204.750 ;
        RECT 110.135 204.280 110.385 204.740 ;
        RECT 110.575 204.490 110.905 204.920 ;
        RECT 111.075 204.950 113.045 205.120 ;
        RECT 111.075 204.450 111.245 204.950 ;
        RECT 111.455 204.280 111.705 204.740 ;
        RECT 111.915 204.450 112.085 204.950 ;
        RECT 112.385 204.280 112.635 204.740 ;
        RECT 112.875 204.450 113.045 204.950 ;
        RECT 113.305 204.450 113.580 205.420 ;
        RECT 113.750 205.250 114.410 205.420 ;
        RECT 114.670 205.300 114.915 205.590 ;
        RECT 114.240 205.130 114.410 205.250 ;
        RECT 115.085 205.130 115.415 205.420 ;
        RECT 113.790 204.280 114.070 205.080 ;
        RECT 114.240 204.960 115.415 205.130 ;
        RECT 115.675 205.030 115.845 205.590 ;
        RECT 114.240 204.460 115.855 204.790 ;
        RECT 116.095 204.280 116.355 205.420 ;
        RECT 116.985 204.280 117.275 205.445 ;
        RECT 117.445 204.280 117.785 205.355 ;
        RECT 117.955 204.995 118.195 205.590 ;
        RECT 118.390 205.130 118.710 205.420 ;
        RECT 118.880 205.300 119.620 205.920 ;
        RECT 119.790 205.590 120.170 205.920 ;
        RECT 120.340 205.590 120.615 205.920 ;
        RECT 120.340 205.420 120.510 205.590 ;
        RECT 120.785 205.420 120.955 206.155 ;
        RECT 119.850 205.250 120.510 205.420 ;
        RECT 119.850 205.130 120.020 205.250 ;
        RECT 118.390 204.960 120.020 205.130 ;
        RECT 117.970 204.500 120.020 204.790 ;
        RECT 120.190 204.280 120.470 205.080 ;
        RECT 120.680 204.450 120.955 205.420 ;
        RECT 121.125 206.155 121.400 206.500 ;
        RECT 121.590 206.430 121.965 206.830 ;
        RECT 122.135 206.260 122.305 206.610 ;
        RECT 122.475 206.430 122.805 206.830 ;
        RECT 122.975 206.260 123.235 206.660 ;
        RECT 121.125 205.420 121.295 206.155 ;
        RECT 121.570 206.090 123.235 206.260 ;
        RECT 121.570 205.920 121.740 206.090 ;
        RECT 123.415 206.010 123.745 206.430 ;
        RECT 123.915 206.010 124.175 206.830 ;
        RECT 124.370 206.075 124.605 206.405 ;
        RECT 124.775 206.090 125.105 206.830 ;
        RECT 125.340 206.450 126.535 206.660 ;
        RECT 123.415 205.920 123.665 206.010 ;
        RECT 121.465 205.590 121.740 205.920 ;
        RECT 121.910 205.590 122.735 205.920 ;
        RECT 122.950 205.590 123.665 205.920 ;
        RECT 123.835 205.590 124.170 205.840 ;
        RECT 121.570 205.420 121.740 205.590 ;
        RECT 121.125 204.450 121.400 205.420 ;
        RECT 121.570 205.250 122.230 205.420 ;
        RECT 122.490 205.300 122.735 205.590 ;
        RECT 122.060 205.130 122.230 205.250 ;
        RECT 122.905 205.130 123.235 205.420 ;
        RECT 121.610 204.280 121.890 205.080 ;
        RECT 122.060 204.960 123.235 205.130 ;
        RECT 123.495 205.030 123.665 205.590 ;
        RECT 124.370 205.420 124.540 206.075 ;
        RECT 125.340 206.010 125.615 206.450 ;
        RECT 125.785 206.010 126.115 206.280 ;
        RECT 126.285 206.220 126.535 206.450 ;
        RECT 126.705 206.390 126.875 206.830 ;
        RECT 127.045 206.220 127.395 206.660 ;
        RECT 126.285 206.010 127.395 206.220 ;
        RECT 127.605 206.010 127.835 206.830 ;
        RECT 128.005 206.030 128.335 206.660 ;
        RECT 125.785 205.980 126.070 206.010 ;
        RECT 124.715 205.590 125.060 205.920 ;
        RECT 125.290 205.420 125.620 205.840 ;
        RECT 122.060 204.460 123.675 204.790 ;
        RECT 123.915 204.280 124.175 205.420 ;
        RECT 124.370 205.250 125.620 205.420 ;
        RECT 124.370 205.055 124.670 205.250 ;
        RECT 125.790 205.080 126.070 205.980 ;
        RECT 126.250 205.640 127.395 205.840 ;
        RECT 126.250 205.260 126.440 205.640 ;
        RECT 127.585 205.590 127.915 205.840 ;
        RECT 128.085 205.430 128.335 206.030 ;
        RECT 128.505 206.010 128.715 206.830 ;
        RECT 128.955 206.020 129.225 206.830 ;
        RECT 129.395 206.020 129.725 206.660 ;
        RECT 129.895 206.020 130.135 206.830 ;
        RECT 130.335 206.020 130.605 206.830 ;
        RECT 130.775 206.020 131.105 206.660 ;
        RECT 131.275 206.020 131.515 206.830 ;
        RECT 132.715 206.280 132.885 206.660 ;
        RECT 133.100 206.450 133.430 206.830 ;
        RECT 132.715 206.110 133.430 206.280 ;
        RECT 128.945 205.590 129.295 205.840 ;
        RECT 126.620 205.080 126.895 205.420 ;
        RECT 124.840 204.280 125.095 205.080 ;
        RECT 125.295 204.910 126.895 205.080 ;
        RECT 125.295 204.450 125.625 204.910 ;
        RECT 125.795 204.280 126.370 204.740 ;
        RECT 126.540 204.450 126.895 204.910 ;
        RECT 127.065 204.280 127.395 205.420 ;
        RECT 127.605 204.280 127.835 205.420 ;
        RECT 128.005 204.450 128.335 205.430 ;
        RECT 129.465 205.420 129.635 206.020 ;
        RECT 129.805 205.590 130.155 205.840 ;
        RECT 130.325 205.590 130.675 205.840 ;
        RECT 130.845 205.420 131.015 206.020 ;
        RECT 131.185 205.590 131.535 205.840 ;
        RECT 132.625 205.560 132.980 205.930 ;
        RECT 133.260 205.920 133.430 206.110 ;
        RECT 133.600 206.085 133.855 206.660 ;
        RECT 133.260 205.590 133.515 205.920 ;
        RECT 128.505 204.280 128.715 205.420 ;
        RECT 128.955 204.280 129.285 205.420 ;
        RECT 129.465 205.250 130.145 205.420 ;
        RECT 129.815 204.465 130.145 205.250 ;
        RECT 130.335 204.280 130.665 205.420 ;
        RECT 130.845 205.250 131.525 205.420 ;
        RECT 133.260 205.380 133.430 205.590 ;
        RECT 131.195 204.465 131.525 205.250 ;
        RECT 132.715 205.210 133.430 205.380 ;
        RECT 133.685 205.355 133.855 206.085 ;
        RECT 134.030 205.990 134.290 206.830 ;
        RECT 134.465 206.090 134.850 206.660 ;
        RECT 135.020 206.370 135.345 206.830 ;
        RECT 135.865 206.200 136.145 206.660 ;
        RECT 132.715 204.450 132.885 205.210 ;
        RECT 133.100 204.280 133.430 205.040 ;
        RECT 133.600 204.450 133.855 205.355 ;
        RECT 134.030 204.280 134.290 205.430 ;
        RECT 134.465 205.420 134.745 206.090 ;
        RECT 135.020 206.030 136.145 206.200 ;
        RECT 135.020 205.920 135.470 206.030 ;
        RECT 134.915 205.590 135.470 205.920 ;
        RECT 136.335 205.860 136.735 206.660 ;
        RECT 137.135 206.370 137.405 206.830 ;
        RECT 137.575 206.200 137.860 206.660 ;
        RECT 134.465 204.450 134.850 205.420 ;
        RECT 135.020 205.130 135.470 205.590 ;
        RECT 135.640 205.300 136.735 205.860 ;
        RECT 135.020 204.910 136.145 205.130 ;
        RECT 135.020 204.280 135.345 204.740 ;
        RECT 135.865 204.450 136.145 204.910 ;
        RECT 136.335 204.450 136.735 205.300 ;
        RECT 136.905 206.030 137.860 206.200 ;
        RECT 138.145 206.060 140.735 206.830 ;
        RECT 140.995 206.280 141.165 206.660 ;
        RECT 141.380 206.450 141.710 206.830 ;
        RECT 140.995 206.110 141.710 206.280 ;
        RECT 136.905 205.130 137.115 206.030 ;
        RECT 137.285 205.300 137.975 205.860 ;
        RECT 138.145 205.540 139.355 206.060 ;
        RECT 139.525 205.370 140.735 205.890 ;
        RECT 140.905 205.560 141.260 205.930 ;
        RECT 141.540 205.920 141.710 206.110 ;
        RECT 141.880 206.085 142.135 206.660 ;
        RECT 141.540 205.590 141.795 205.920 ;
        RECT 141.540 205.380 141.710 205.590 ;
        RECT 136.905 204.910 137.860 205.130 ;
        RECT 137.135 204.280 137.405 204.740 ;
        RECT 137.575 204.450 137.860 204.910 ;
        RECT 138.145 204.280 140.735 205.370 ;
        RECT 140.995 205.210 141.710 205.380 ;
        RECT 141.965 205.355 142.135 206.085 ;
        RECT 142.310 205.990 142.570 206.830 ;
        RECT 142.745 206.105 143.035 206.830 ;
        RECT 143.205 206.080 144.415 206.830 ;
        RECT 144.675 206.280 144.845 206.660 ;
        RECT 145.060 206.450 145.390 206.830 ;
        RECT 144.675 206.110 145.390 206.280 ;
        RECT 143.205 205.540 143.725 206.080 ;
        RECT 140.995 204.450 141.165 205.210 ;
        RECT 141.380 204.280 141.710 205.040 ;
        RECT 141.880 204.450 142.135 205.355 ;
        RECT 142.310 204.280 142.570 205.430 ;
        RECT 142.745 204.280 143.035 205.445 ;
        RECT 143.895 205.370 144.415 205.910 ;
        RECT 144.585 205.560 144.940 205.930 ;
        RECT 145.220 205.920 145.390 206.110 ;
        RECT 145.560 206.085 145.815 206.660 ;
        RECT 145.220 205.590 145.475 205.920 ;
        RECT 145.220 205.380 145.390 205.590 ;
        RECT 143.205 204.280 144.415 205.370 ;
        RECT 144.675 205.210 145.390 205.380 ;
        RECT 145.645 205.355 145.815 206.085 ;
        RECT 145.990 205.990 146.250 206.830 ;
        RECT 146.425 206.080 147.635 206.830 ;
        RECT 144.675 204.450 144.845 205.210 ;
        RECT 145.060 204.280 145.390 205.040 ;
        RECT 145.560 204.450 145.815 205.355 ;
        RECT 145.990 204.280 146.250 205.430 ;
        RECT 146.425 205.370 146.945 205.910 ;
        RECT 147.115 205.540 147.635 206.080 ;
        RECT 146.425 204.280 147.635 205.370 ;
        RECT 13.860 204.110 147.720 204.280 ;
        RECT 13.945 203.020 15.155 204.110 ;
        RECT 13.945 202.310 14.465 202.850 ;
        RECT 14.635 202.480 15.155 203.020 ;
        RECT 15.330 202.960 15.590 204.110 ;
        RECT 15.765 203.035 16.020 203.940 ;
        RECT 16.190 203.350 16.520 204.110 ;
        RECT 16.735 203.180 16.905 203.940 ;
        RECT 17.630 203.440 17.885 203.940 ;
        RECT 18.055 203.610 18.385 204.110 ;
        RECT 17.630 203.270 18.380 203.440 ;
        RECT 13.945 201.560 15.155 202.310 ;
        RECT 15.330 201.560 15.590 202.400 ;
        RECT 15.765 202.305 15.935 203.035 ;
        RECT 16.190 203.010 16.905 203.180 ;
        RECT 16.190 202.800 16.360 203.010 ;
        RECT 16.105 202.470 16.360 202.800 ;
        RECT 15.765 201.730 16.020 202.305 ;
        RECT 16.190 202.280 16.360 202.470 ;
        RECT 16.640 202.460 16.995 202.830 ;
        RECT 17.630 202.450 17.980 203.100 ;
        RECT 18.150 202.280 18.380 203.270 ;
        RECT 16.190 202.110 16.905 202.280 ;
        RECT 16.190 201.560 16.520 201.940 ;
        RECT 16.735 201.730 16.905 202.110 ;
        RECT 17.630 202.110 18.380 202.280 ;
        RECT 17.630 201.820 17.885 202.110 ;
        RECT 18.055 201.560 18.385 201.940 ;
        RECT 18.555 201.820 18.725 203.940 ;
        RECT 18.895 203.140 19.220 203.925 ;
        RECT 19.390 203.650 19.640 204.110 ;
        RECT 19.810 203.610 20.060 203.940 ;
        RECT 20.275 203.610 20.955 203.940 ;
        RECT 19.810 203.480 19.980 203.610 ;
        RECT 19.585 203.310 19.980 203.480 ;
        RECT 18.955 202.090 19.415 203.140 ;
        RECT 19.585 201.950 19.755 203.310 ;
        RECT 20.150 203.050 20.615 203.440 ;
        RECT 19.925 202.240 20.275 202.860 ;
        RECT 20.445 202.460 20.615 203.050 ;
        RECT 20.785 202.830 20.955 203.610 ;
        RECT 21.125 203.510 21.295 203.850 ;
        RECT 21.530 203.680 21.860 204.110 ;
        RECT 22.030 203.510 22.200 203.850 ;
        RECT 22.495 203.650 22.865 204.110 ;
        RECT 21.125 203.340 22.200 203.510 ;
        RECT 23.035 203.480 23.205 203.940 ;
        RECT 23.440 203.600 24.310 203.940 ;
        RECT 24.480 203.650 24.730 204.110 ;
        RECT 22.645 203.310 23.205 203.480 ;
        RECT 22.645 203.170 22.815 203.310 ;
        RECT 21.315 203.000 22.815 203.170 ;
        RECT 23.510 203.140 23.970 203.430 ;
        RECT 20.785 202.660 22.475 202.830 ;
        RECT 20.445 202.240 20.800 202.460 ;
        RECT 20.970 201.950 21.140 202.660 ;
        RECT 21.345 202.240 22.135 202.490 ;
        RECT 22.305 202.480 22.475 202.660 ;
        RECT 22.645 202.310 22.815 203.000 ;
        RECT 19.085 201.560 19.415 201.920 ;
        RECT 19.585 201.780 20.080 201.950 ;
        RECT 20.285 201.780 21.140 201.950 ;
        RECT 22.015 201.560 22.345 202.020 ;
        RECT 22.555 201.920 22.815 202.310 ;
        RECT 23.005 203.130 23.970 203.140 ;
        RECT 24.140 203.220 24.310 203.600 ;
        RECT 24.900 203.560 25.070 203.850 ;
        RECT 25.250 203.730 25.580 204.110 ;
        RECT 24.900 203.390 25.700 203.560 ;
        RECT 23.005 202.970 23.680 203.130 ;
        RECT 24.140 203.050 25.360 203.220 ;
        RECT 23.005 202.180 23.215 202.970 ;
        RECT 24.140 202.960 24.310 203.050 ;
        RECT 23.385 202.180 23.735 202.800 ;
        RECT 23.905 202.790 24.310 202.960 ;
        RECT 23.905 202.010 24.075 202.790 ;
        RECT 24.245 202.340 24.465 202.620 ;
        RECT 24.645 202.510 25.185 202.880 ;
        RECT 25.530 202.800 25.700 203.390 ;
        RECT 25.920 202.970 26.225 204.110 ;
        RECT 26.395 202.920 26.650 203.800 ;
        RECT 26.825 202.945 27.115 204.110 ;
        RECT 27.290 202.970 27.625 203.940 ;
        RECT 27.795 202.970 27.965 204.110 ;
        RECT 28.135 203.770 30.165 203.940 ;
        RECT 25.530 202.770 26.270 202.800 ;
        RECT 24.245 202.170 24.775 202.340 ;
        RECT 22.555 201.750 22.905 201.920 ;
        RECT 23.125 201.730 24.075 202.010 ;
        RECT 24.245 201.560 24.435 202.000 ;
        RECT 24.605 201.940 24.775 202.170 ;
        RECT 24.945 202.110 25.185 202.510 ;
        RECT 25.355 202.470 26.270 202.770 ;
        RECT 25.355 202.295 25.680 202.470 ;
        RECT 25.355 201.940 25.675 202.295 ;
        RECT 26.440 202.270 26.650 202.920 ;
        RECT 27.290 202.300 27.460 202.970 ;
        RECT 28.135 202.800 28.305 203.770 ;
        RECT 27.630 202.470 27.885 202.800 ;
        RECT 28.110 202.470 28.305 202.800 ;
        RECT 28.475 203.430 29.600 203.600 ;
        RECT 27.715 202.300 27.885 202.470 ;
        RECT 28.475 202.300 28.645 203.430 ;
        RECT 24.605 201.770 25.675 201.940 ;
        RECT 25.920 201.560 26.225 202.020 ;
        RECT 26.395 201.740 26.650 202.270 ;
        RECT 26.825 201.560 27.115 202.285 ;
        RECT 27.290 201.730 27.545 202.300 ;
        RECT 27.715 202.130 28.645 202.300 ;
        RECT 28.815 203.090 29.825 203.260 ;
        RECT 28.815 202.290 28.985 203.090 ;
        RECT 29.190 202.750 29.465 202.890 ;
        RECT 29.185 202.580 29.465 202.750 ;
        RECT 28.470 202.095 28.645 202.130 ;
        RECT 27.715 201.560 28.045 201.960 ;
        RECT 28.470 201.730 29.000 202.095 ;
        RECT 29.190 201.730 29.465 202.580 ;
        RECT 29.635 201.730 29.825 203.090 ;
        RECT 29.995 203.105 30.165 203.770 ;
        RECT 30.335 203.350 30.505 204.110 ;
        RECT 30.740 203.350 31.255 203.760 ;
        RECT 29.995 202.915 30.745 203.105 ;
        RECT 30.915 202.540 31.255 203.350 ;
        RECT 30.025 202.370 31.255 202.540 ;
        RECT 31.425 203.520 32.125 203.940 ;
        RECT 32.325 203.750 32.655 204.110 ;
        RECT 32.825 203.520 33.155 203.920 ;
        RECT 31.425 203.290 33.155 203.520 ;
        RECT 30.005 201.560 30.515 202.095 ;
        RECT 30.735 201.765 30.980 202.370 ;
        RECT 31.425 202.320 31.630 203.290 ;
        RECT 31.800 202.550 32.130 203.090 ;
        RECT 32.305 202.800 32.630 203.090 ;
        RECT 32.825 203.070 33.155 203.290 ;
        RECT 33.325 202.800 33.495 203.725 ;
        RECT 33.675 203.050 34.005 204.110 ;
        RECT 34.275 203.365 34.545 204.110 ;
        RECT 35.175 204.105 41.450 204.110 ;
        RECT 34.715 203.195 35.005 203.935 ;
        RECT 35.175 203.380 35.430 204.105 ;
        RECT 35.615 203.210 35.875 203.935 ;
        RECT 36.045 203.380 36.290 204.105 ;
        RECT 36.475 203.210 36.735 203.935 ;
        RECT 36.905 203.380 37.150 204.105 ;
        RECT 37.335 203.210 37.595 203.935 ;
        RECT 37.765 203.380 38.010 204.105 ;
        RECT 38.180 203.210 38.440 203.935 ;
        RECT 38.610 203.380 38.870 204.105 ;
        RECT 39.040 203.210 39.300 203.935 ;
        RECT 39.470 203.380 39.730 204.105 ;
        RECT 39.900 203.210 40.160 203.935 ;
        RECT 40.330 203.380 40.590 204.105 ;
        RECT 40.760 203.210 41.020 203.935 ;
        RECT 41.190 203.310 41.450 204.105 ;
        RECT 35.615 203.195 41.020 203.210 ;
        RECT 34.275 202.970 41.020 203.195 ;
        RECT 32.305 202.470 32.800 202.800 ;
        RECT 33.120 202.470 33.495 202.800 ;
        RECT 33.705 202.470 34.015 202.800 ;
        RECT 34.275 202.380 35.440 202.970 ;
        RECT 41.620 202.800 41.870 203.935 ;
        RECT 42.050 203.300 42.310 204.110 ;
        RECT 42.485 202.800 42.730 203.940 ;
        RECT 42.910 203.300 43.205 204.110 ;
        RECT 43.440 203.240 43.725 204.110 ;
        RECT 43.895 203.480 44.155 203.940 ;
        RECT 44.330 203.650 44.585 204.110 ;
        RECT 44.755 203.480 45.015 203.940 ;
        RECT 43.895 203.310 45.015 203.480 ;
        RECT 45.185 203.310 45.495 204.110 ;
        RECT 43.895 203.060 44.155 203.310 ;
        RECT 45.665 203.140 45.975 203.940 ;
        RECT 43.400 202.890 44.155 203.060 ;
        RECT 44.945 202.970 45.975 203.140 ;
        RECT 46.605 202.970 46.865 204.110 ;
        RECT 47.035 203.140 47.365 203.940 ;
        RECT 47.535 203.310 47.705 204.110 ;
        RECT 47.875 203.140 48.205 203.940 ;
        RECT 48.375 203.310 48.630 204.110 ;
        RECT 47.035 202.970 48.735 203.140 ;
        RECT 48.965 202.970 49.175 204.110 ;
        RECT 35.610 202.550 42.730 202.800 ;
        RECT 31.425 201.730 32.135 202.320 ;
        RECT 32.645 202.090 34.005 202.300 ;
        RECT 34.275 202.210 41.020 202.380 ;
        RECT 32.645 201.730 32.975 202.090 ;
        RECT 33.175 201.560 33.505 201.920 ;
        RECT 33.675 201.730 34.005 202.090 ;
        RECT 34.275 201.560 34.575 202.040 ;
        RECT 34.745 201.755 35.005 202.210 ;
        RECT 35.175 201.560 35.435 202.040 ;
        RECT 35.615 201.755 35.875 202.210 ;
        RECT 36.045 201.560 36.295 202.040 ;
        RECT 36.475 201.755 36.735 202.210 ;
        RECT 36.905 201.560 37.155 202.040 ;
        RECT 37.335 201.755 37.595 202.210 ;
        RECT 37.765 201.560 38.010 202.040 ;
        RECT 38.180 201.755 38.455 202.210 ;
        RECT 38.625 201.560 38.870 202.040 ;
        RECT 39.040 201.755 39.300 202.210 ;
        RECT 39.470 201.560 39.730 202.040 ;
        RECT 39.900 201.755 40.160 202.210 ;
        RECT 40.330 201.560 40.590 202.040 ;
        RECT 40.760 201.755 41.020 202.210 ;
        RECT 41.190 201.560 41.450 202.120 ;
        RECT 41.620 201.740 41.870 202.550 ;
        RECT 42.050 201.560 42.310 202.085 ;
        RECT 42.480 201.740 42.730 202.550 ;
        RECT 42.900 202.240 43.215 202.800 ;
        RECT 43.400 202.380 43.805 202.890 ;
        RECT 44.945 202.720 45.115 202.970 ;
        RECT 43.975 202.550 45.115 202.720 ;
        RECT 43.400 202.210 45.050 202.380 ;
        RECT 45.285 202.230 45.635 202.800 ;
        RECT 42.910 201.560 43.215 202.070 ;
        RECT 43.445 201.560 43.725 202.040 ;
        RECT 43.895 201.820 44.155 202.210 ;
        RECT 44.330 201.560 44.585 202.040 ;
        RECT 44.755 201.820 45.050 202.210 ;
        RECT 45.805 202.060 45.975 202.970 ;
        RECT 46.605 202.550 47.365 202.800 ;
        RECT 47.535 202.550 48.285 202.800 ;
        RECT 48.455 202.380 48.735 202.970 ;
        RECT 49.345 202.960 49.675 203.940 ;
        RECT 49.845 202.970 50.075 204.110 ;
        RECT 50.295 203.140 50.625 203.925 ;
        RECT 50.295 202.970 50.975 203.140 ;
        RECT 51.155 202.970 51.485 204.110 ;
        RECT 45.230 201.560 45.505 202.040 ;
        RECT 45.675 201.730 45.975 202.060 ;
        RECT 46.605 202.190 47.705 202.360 ;
        RECT 46.605 201.730 46.945 202.190 ;
        RECT 47.115 201.560 47.285 202.020 ;
        RECT 47.455 201.940 47.705 202.190 ;
        RECT 47.875 202.130 48.735 202.380 ;
        RECT 48.295 201.940 48.625 201.960 ;
        RECT 47.455 201.730 48.625 201.940 ;
        RECT 48.965 201.560 49.175 202.380 ;
        RECT 49.345 202.360 49.595 202.960 ;
        RECT 49.765 202.550 50.095 202.800 ;
        RECT 50.285 202.550 50.635 202.800 ;
        RECT 49.345 201.730 49.675 202.360 ;
        RECT 49.845 201.560 50.075 202.380 ;
        RECT 50.805 202.370 50.975 202.970 ;
        RECT 52.585 202.945 52.875 204.110 ;
        RECT 53.505 203.140 53.775 203.910 ;
        RECT 53.945 203.330 54.275 204.110 ;
        RECT 54.480 203.505 54.665 203.910 ;
        RECT 54.835 203.685 55.170 204.110 ;
        RECT 54.480 203.330 55.145 203.505 ;
        RECT 53.505 202.970 54.635 203.140 ;
        RECT 51.145 202.550 51.495 202.800 ;
        RECT 50.305 201.560 50.545 202.370 ;
        RECT 50.715 201.730 51.045 202.370 ;
        RECT 51.215 201.560 51.485 202.370 ;
        RECT 52.585 201.560 52.875 202.285 ;
        RECT 53.505 202.060 53.675 202.970 ;
        RECT 53.845 202.220 54.205 202.800 ;
        RECT 54.385 202.470 54.635 202.970 ;
        RECT 54.805 202.300 55.145 203.330 ;
        RECT 55.350 203.310 55.665 204.110 ;
        RECT 55.930 203.755 57.010 203.925 ;
        RECT 55.930 203.140 56.100 203.755 ;
        RECT 54.460 202.130 55.145 202.300 ;
        RECT 55.345 202.130 55.615 203.140 ;
        RECT 55.785 202.970 56.100 203.140 ;
        RECT 55.785 202.300 55.955 202.970 ;
        RECT 56.270 202.800 56.505 203.480 ;
        RECT 56.675 202.970 57.010 203.755 ;
        RECT 57.390 203.140 57.720 203.940 ;
        RECT 57.890 203.310 58.220 204.110 ;
        RECT 58.520 203.140 58.850 203.940 ;
        RECT 59.495 203.310 59.745 204.110 ;
        RECT 57.390 202.970 59.825 203.140 ;
        RECT 60.015 202.970 60.185 204.110 ;
        RECT 60.355 202.970 60.695 203.940 ;
        RECT 60.875 203.300 61.170 204.110 ;
        RECT 56.125 202.470 56.505 202.800 ;
        RECT 56.675 202.470 57.010 202.800 ;
        RECT 57.185 202.550 57.535 202.800 ;
        RECT 57.720 202.340 57.890 202.970 ;
        RECT 58.060 202.550 58.390 202.750 ;
        RECT 58.560 202.550 58.890 202.750 ;
        RECT 59.060 202.550 59.480 202.750 ;
        RECT 59.655 202.720 59.825 202.970 ;
        RECT 59.655 202.550 60.350 202.720 ;
        RECT 55.785 202.130 57.010 202.300 ;
        RECT 53.505 201.730 53.765 202.060 ;
        RECT 53.975 201.560 54.250 202.040 ;
        RECT 54.460 201.730 54.665 202.130 ;
        RECT 54.835 201.560 55.170 201.960 ;
        RECT 55.415 201.560 55.745 201.960 ;
        RECT 55.915 201.860 56.085 202.130 ;
        RECT 56.255 201.560 56.585 201.960 ;
        RECT 56.755 201.860 57.010 202.130 ;
        RECT 57.390 201.730 57.890 202.340 ;
        RECT 58.520 202.210 59.745 202.380 ;
        RECT 60.520 202.360 60.695 202.970 ;
        RECT 61.350 202.800 61.595 203.940 ;
        RECT 61.770 203.300 62.030 204.110 ;
        RECT 62.630 204.105 68.905 204.110 ;
        RECT 62.210 202.800 62.460 203.935 ;
        RECT 62.630 203.310 62.890 204.105 ;
        RECT 63.060 203.210 63.320 203.935 ;
        RECT 63.490 203.380 63.750 204.105 ;
        RECT 63.920 203.210 64.180 203.935 ;
        RECT 64.350 203.380 64.610 204.105 ;
        RECT 64.780 203.210 65.040 203.935 ;
        RECT 65.210 203.380 65.470 204.105 ;
        RECT 65.640 203.210 65.900 203.935 ;
        RECT 66.070 203.380 66.315 204.105 ;
        RECT 66.485 203.210 66.745 203.935 ;
        RECT 66.930 203.380 67.175 204.105 ;
        RECT 67.345 203.210 67.605 203.935 ;
        RECT 67.790 203.380 68.035 204.105 ;
        RECT 68.205 203.210 68.465 203.935 ;
        RECT 68.650 203.380 68.905 204.105 ;
        RECT 63.060 203.195 68.465 203.210 ;
        RECT 69.075 203.195 69.365 203.935 ;
        RECT 69.535 203.365 69.805 204.110 ;
        RECT 63.060 202.970 69.805 203.195 ;
        RECT 58.520 201.730 58.850 202.210 ;
        RECT 59.020 201.560 59.245 202.020 ;
        RECT 59.415 201.730 59.745 202.210 ;
        RECT 59.935 201.560 60.185 202.360 ;
        RECT 60.355 201.730 60.695 202.360 ;
        RECT 60.865 202.240 61.180 202.800 ;
        RECT 61.350 202.550 68.470 202.800 ;
        RECT 60.865 201.560 61.170 202.070 ;
        RECT 61.350 201.740 61.600 202.550 ;
        RECT 61.770 201.560 62.030 202.085 ;
        RECT 62.210 201.740 62.460 202.550 ;
        RECT 68.640 202.380 69.805 202.970 ;
        RECT 63.060 202.210 69.805 202.380 ;
        RECT 70.065 202.970 70.340 203.940 ;
        RECT 70.550 203.310 70.830 204.110 ;
        RECT 71.000 203.600 72.615 203.930 ;
        RECT 71.000 203.260 72.175 203.430 ;
        RECT 71.000 203.140 71.170 203.260 ;
        RECT 70.510 202.970 71.170 203.140 ;
        RECT 70.065 202.235 70.235 202.970 ;
        RECT 70.510 202.800 70.680 202.970 ;
        RECT 71.430 202.800 71.675 203.090 ;
        RECT 71.845 202.970 72.175 203.260 ;
        RECT 72.435 202.800 72.605 203.360 ;
        RECT 72.855 202.970 73.115 204.110 ;
        RECT 73.285 203.600 74.475 203.890 ;
        RECT 73.305 203.260 74.475 203.430 ;
        RECT 74.645 203.310 74.925 204.110 ;
        RECT 73.305 202.970 73.630 203.260 ;
        RECT 74.305 203.140 74.475 203.260 ;
        RECT 73.800 202.800 73.995 203.090 ;
        RECT 74.305 202.970 74.965 203.140 ;
        RECT 75.135 202.970 75.410 203.940 ;
        RECT 75.590 202.970 75.910 204.110 ;
        RECT 74.795 202.800 74.965 202.970 ;
        RECT 70.405 202.470 70.680 202.800 ;
        RECT 70.850 202.470 71.675 202.800 ;
        RECT 71.890 202.470 72.605 202.800 ;
        RECT 72.775 202.550 73.110 202.800 ;
        RECT 73.285 202.470 73.630 202.800 ;
        RECT 73.800 202.470 74.625 202.800 ;
        RECT 74.795 202.470 75.070 202.800 ;
        RECT 70.510 202.300 70.680 202.470 ;
        RECT 72.355 202.380 72.605 202.470 ;
        RECT 62.630 201.560 62.890 202.120 ;
        RECT 63.060 201.755 63.320 202.210 ;
        RECT 63.490 201.560 63.750 202.040 ;
        RECT 63.920 201.755 64.180 202.210 ;
        RECT 64.350 201.560 64.610 202.040 ;
        RECT 64.780 201.755 65.040 202.210 ;
        RECT 65.210 201.560 65.455 202.040 ;
        RECT 65.625 201.755 65.900 202.210 ;
        RECT 66.070 201.560 66.315 202.040 ;
        RECT 66.485 201.755 66.745 202.210 ;
        RECT 66.925 201.560 67.175 202.040 ;
        RECT 67.345 201.755 67.605 202.210 ;
        RECT 67.785 201.560 68.035 202.040 ;
        RECT 68.205 201.755 68.465 202.210 ;
        RECT 68.645 201.560 68.905 202.040 ;
        RECT 69.075 201.755 69.335 202.210 ;
        RECT 69.505 201.560 69.805 202.040 ;
        RECT 70.065 201.890 70.340 202.235 ;
        RECT 70.510 202.130 72.175 202.300 ;
        RECT 70.530 201.560 70.905 201.960 ;
        RECT 71.075 201.780 71.245 202.130 ;
        RECT 71.415 201.560 71.745 201.960 ;
        RECT 71.915 201.730 72.175 202.130 ;
        RECT 72.355 201.960 72.685 202.380 ;
        RECT 72.855 201.560 73.115 202.380 ;
        RECT 74.795 202.300 74.965 202.470 ;
        RECT 73.300 202.130 74.965 202.300 ;
        RECT 75.240 202.235 75.410 202.970 ;
        RECT 76.090 202.800 76.285 203.850 ;
        RECT 76.465 203.260 76.795 203.940 ;
        RECT 76.995 203.310 77.250 204.110 ;
        RECT 76.465 202.980 76.815 203.260 ;
        RECT 75.650 202.750 75.910 202.800 ;
        RECT 75.645 202.580 75.910 202.750 ;
        RECT 75.650 202.470 75.910 202.580 ;
        RECT 76.090 202.470 76.475 202.800 ;
        RECT 76.645 202.600 76.815 202.980 ;
        RECT 77.005 202.770 77.250 203.130 ;
        RECT 78.345 202.945 78.635 204.110 ;
        RECT 78.805 203.515 79.240 203.940 ;
        RECT 79.410 203.685 79.795 204.110 ;
        RECT 78.805 203.345 79.795 203.515 ;
        RECT 76.645 202.430 77.165 202.600 ;
        RECT 78.805 202.470 79.290 203.175 ;
        RECT 79.460 202.800 79.795 203.345 ;
        RECT 79.965 203.150 80.390 203.940 ;
        RECT 80.560 203.515 80.835 203.940 ;
        RECT 81.005 203.685 81.390 204.110 ;
        RECT 80.560 203.320 81.390 203.515 ;
        RECT 79.965 202.970 80.870 203.150 ;
        RECT 79.460 202.470 79.870 202.800 ;
        RECT 80.040 202.470 80.870 202.970 ;
        RECT 81.040 202.800 81.390 203.320 ;
        RECT 81.560 203.150 81.805 203.940 ;
        RECT 81.995 203.515 82.250 203.940 ;
        RECT 82.420 203.685 82.805 204.110 ;
        RECT 81.995 203.320 82.805 203.515 ;
        RECT 81.560 202.970 82.285 203.150 ;
        RECT 81.040 202.470 81.465 202.800 ;
        RECT 81.635 202.470 82.285 202.970 ;
        RECT 82.455 202.800 82.805 203.320 ;
        RECT 82.975 202.970 83.235 203.940 ;
        RECT 83.405 202.970 83.685 204.110 ;
        RECT 82.455 202.470 82.880 202.800 ;
        RECT 73.300 201.780 73.555 202.130 ;
        RECT 73.725 201.560 74.055 201.960 ;
        RECT 74.225 201.780 74.395 202.130 ;
        RECT 74.565 201.560 74.945 201.960 ;
        RECT 75.135 201.890 75.410 202.235 ;
        RECT 75.590 202.090 76.805 202.260 ;
        RECT 75.590 201.740 75.880 202.090 ;
        RECT 76.075 201.560 76.405 201.920 ;
        RECT 76.575 201.785 76.805 202.090 ;
        RECT 76.995 202.070 77.165 202.430 ;
        RECT 79.460 202.300 79.795 202.470 ;
        RECT 80.040 202.300 80.390 202.470 ;
        RECT 81.040 202.300 81.390 202.470 ;
        RECT 81.635 202.300 81.805 202.470 ;
        RECT 82.455 202.300 82.805 202.470 ;
        RECT 83.050 202.300 83.235 202.970 ;
        RECT 83.855 202.960 84.185 203.940 ;
        RECT 84.355 202.970 84.615 204.110 ;
        RECT 84.845 202.970 85.055 204.110 ;
        RECT 85.225 202.960 85.555 203.940 ;
        RECT 85.725 202.970 85.955 204.110 ;
        RECT 87.090 203.310 87.345 204.110 ;
        RECT 87.545 203.260 87.875 203.940 ;
        RECT 83.920 202.920 84.095 202.960 ;
        RECT 83.415 202.530 83.750 202.800 ;
        RECT 83.920 202.360 84.090 202.920 ;
        RECT 84.260 202.550 84.595 202.800 ;
        RECT 76.995 201.900 77.195 202.070 ;
        RECT 76.995 201.865 77.165 201.900 ;
        RECT 78.345 201.560 78.635 202.285 ;
        RECT 78.805 202.130 79.795 202.300 ;
        RECT 78.805 201.730 79.240 202.130 ;
        RECT 79.410 201.560 79.795 201.960 ;
        RECT 79.965 201.730 80.390 202.300 ;
        RECT 80.580 202.130 81.390 202.300 ;
        RECT 80.580 201.730 80.835 202.130 ;
        RECT 81.005 201.560 81.390 201.960 ;
        RECT 81.560 201.730 81.805 202.300 ;
        RECT 81.995 202.130 82.805 202.300 ;
        RECT 81.995 201.730 82.250 202.130 ;
        RECT 82.420 201.560 82.805 201.960 ;
        RECT 82.975 201.730 83.235 202.300 ;
        RECT 83.405 201.560 83.715 202.360 ;
        RECT 83.920 201.730 84.615 202.360 ;
        RECT 84.845 201.560 85.055 202.380 ;
        RECT 85.225 202.360 85.475 202.960 ;
        RECT 85.645 202.550 85.975 202.800 ;
        RECT 87.090 202.770 87.335 203.130 ;
        RECT 87.525 202.980 87.875 203.260 ;
        RECT 87.525 202.600 87.695 202.980 ;
        RECT 88.055 202.800 88.250 203.850 ;
        RECT 88.430 202.970 88.750 204.110 ;
        RECT 88.925 202.970 89.185 204.110 ;
        RECT 89.355 202.960 89.685 203.940 ;
        RECT 89.855 202.970 90.135 204.110 ;
        RECT 90.305 202.970 90.585 204.110 ;
        RECT 90.755 202.960 91.085 203.940 ;
        RECT 91.255 202.970 91.515 204.110 ;
        RECT 92.145 202.970 92.405 204.110 ;
        RECT 92.575 202.960 92.905 203.940 ;
        RECT 93.075 202.970 93.355 204.110 ;
        RECT 93.525 202.970 93.785 204.110 ;
        RECT 93.955 202.960 94.285 203.940 ;
        RECT 94.455 202.970 94.735 204.110 ;
        RECT 94.910 203.160 95.175 203.930 ;
        RECT 95.345 203.390 95.675 204.110 ;
        RECT 95.865 203.570 96.125 203.930 ;
        RECT 96.295 203.740 96.625 204.110 ;
        RECT 96.795 203.570 97.055 203.930 ;
        RECT 95.865 203.340 97.055 203.570 ;
        RECT 97.625 203.160 97.915 203.930 ;
        RECT 87.175 202.430 87.695 202.600 ;
        RECT 87.865 202.470 88.250 202.800 ;
        RECT 88.430 202.750 88.690 202.800 ;
        RECT 88.430 202.580 88.695 202.750 ;
        RECT 88.430 202.470 88.690 202.580 ;
        RECT 88.945 202.550 89.280 202.800 ;
        RECT 85.225 201.730 85.555 202.360 ;
        RECT 85.725 201.560 85.955 202.380 ;
        RECT 87.175 201.865 87.345 202.430 ;
        RECT 89.450 202.360 89.620 202.960 ;
        RECT 89.790 202.530 90.125 202.800 ;
        RECT 90.315 202.530 90.650 202.800 ;
        RECT 90.820 202.360 90.990 202.960 ;
        RECT 91.160 202.550 91.495 202.800 ;
        RECT 92.165 202.550 92.500 202.800 ;
        RECT 92.670 202.360 92.840 202.960 ;
        RECT 93.010 202.530 93.345 202.800 ;
        RECT 93.545 202.550 93.880 202.800 ;
        RECT 94.050 202.360 94.220 202.960 ;
        RECT 94.390 202.530 94.725 202.800 ;
        RECT 87.535 202.090 88.750 202.260 ;
        RECT 87.535 201.785 87.765 202.090 ;
        RECT 87.935 201.560 88.265 201.920 ;
        RECT 88.460 201.740 88.750 202.090 ;
        RECT 88.925 201.730 89.620 202.360 ;
        RECT 89.825 201.560 90.135 202.360 ;
        RECT 90.305 201.560 90.615 202.360 ;
        RECT 90.820 201.730 91.515 202.360 ;
        RECT 92.145 201.730 92.840 202.360 ;
        RECT 93.045 201.560 93.355 202.360 ;
        RECT 93.525 201.730 94.220 202.360 ;
        RECT 94.425 201.560 94.735 202.360 ;
        RECT 94.910 201.740 95.245 203.160 ;
        RECT 95.420 202.980 97.915 203.160 ;
        RECT 98.130 203.160 98.395 203.930 ;
        RECT 98.565 203.390 98.895 204.110 ;
        RECT 99.085 203.570 99.345 203.930 ;
        RECT 99.515 203.740 99.845 204.110 ;
        RECT 100.015 203.570 100.275 203.930 ;
        RECT 99.085 203.340 100.275 203.570 ;
        RECT 100.845 203.160 101.135 203.930 ;
        RECT 95.420 202.290 95.645 202.980 ;
        RECT 95.845 202.470 96.125 202.800 ;
        RECT 96.305 202.470 96.880 202.800 ;
        RECT 97.060 202.470 97.495 202.800 ;
        RECT 97.675 202.470 97.945 202.800 ;
        RECT 95.420 202.100 97.905 202.290 ;
        RECT 95.425 201.560 96.170 201.930 ;
        RECT 96.735 201.740 96.990 202.100 ;
        RECT 97.170 201.560 97.500 201.930 ;
        RECT 97.680 201.740 97.905 202.100 ;
        RECT 98.130 201.740 98.465 203.160 ;
        RECT 98.640 202.980 101.135 203.160 ;
        RECT 98.640 202.290 98.865 202.980 ;
        RECT 102.265 202.970 102.545 204.110 ;
        RECT 102.715 202.960 103.045 203.940 ;
        RECT 103.215 202.970 103.475 204.110 ;
        RECT 99.065 202.470 99.345 202.800 ;
        RECT 99.525 202.470 100.100 202.800 ;
        RECT 100.280 202.470 100.715 202.800 ;
        RECT 100.895 202.470 101.165 202.800 ;
        RECT 102.275 202.530 102.610 202.800 ;
        RECT 102.780 202.360 102.950 202.960 ;
        RECT 104.105 202.945 104.395 204.110 ;
        RECT 104.570 202.970 104.905 203.940 ;
        RECT 105.075 202.970 105.245 204.110 ;
        RECT 105.415 203.770 107.445 203.940 ;
        RECT 103.120 202.550 103.455 202.800 ;
        RECT 98.640 202.100 101.125 202.290 ;
        RECT 98.645 201.560 99.390 201.930 ;
        RECT 99.955 201.740 100.210 202.100 ;
        RECT 100.390 201.560 100.720 201.930 ;
        RECT 100.900 201.740 101.125 202.100 ;
        RECT 102.265 201.560 102.575 202.360 ;
        RECT 102.780 201.730 103.475 202.360 ;
        RECT 104.570 202.300 104.740 202.970 ;
        RECT 105.415 202.800 105.585 203.770 ;
        RECT 104.910 202.470 105.165 202.800 ;
        RECT 105.390 202.470 105.585 202.800 ;
        RECT 105.755 203.430 106.880 203.600 ;
        RECT 104.995 202.300 105.165 202.470 ;
        RECT 105.755 202.300 105.925 203.430 ;
        RECT 104.105 201.560 104.395 202.285 ;
        RECT 104.570 201.730 104.825 202.300 ;
        RECT 104.995 202.130 105.925 202.300 ;
        RECT 106.095 203.090 107.105 203.260 ;
        RECT 106.095 202.290 106.265 203.090 ;
        RECT 106.470 202.410 106.745 202.890 ;
        RECT 106.465 202.240 106.745 202.410 ;
        RECT 105.750 202.095 105.925 202.130 ;
        RECT 104.995 201.560 105.325 201.960 ;
        RECT 105.750 201.730 106.280 202.095 ;
        RECT 106.470 201.730 106.745 202.240 ;
        RECT 106.915 201.730 107.105 203.090 ;
        RECT 107.275 203.105 107.445 203.770 ;
        RECT 107.615 203.350 107.785 204.110 ;
        RECT 108.020 203.350 108.535 203.760 ;
        RECT 107.275 202.915 108.025 203.105 ;
        RECT 108.195 202.540 108.535 203.350 ;
        RECT 108.765 202.970 108.975 204.110 ;
        RECT 107.305 202.370 108.535 202.540 ;
        RECT 109.145 202.960 109.475 203.940 ;
        RECT 109.645 202.970 109.875 204.110 ;
        RECT 110.095 203.050 110.425 203.900 ;
        RECT 107.285 201.560 107.795 202.095 ;
        RECT 108.015 201.765 108.260 202.370 ;
        RECT 108.765 201.560 108.975 202.380 ;
        RECT 109.145 202.360 109.395 202.960 ;
        RECT 109.565 202.550 109.895 202.800 ;
        RECT 109.145 201.730 109.475 202.360 ;
        RECT 109.645 201.560 109.875 202.380 ;
        RECT 110.095 202.285 110.285 203.050 ;
        RECT 110.595 202.970 110.845 204.110 ;
        RECT 111.035 203.470 111.285 203.890 ;
        RECT 111.515 203.640 111.845 204.110 ;
        RECT 112.075 203.470 112.325 203.890 ;
        RECT 111.035 203.300 112.325 203.470 ;
        RECT 112.505 203.470 112.835 203.900 ;
        RECT 112.505 203.300 112.960 203.470 ;
        RECT 111.025 202.800 111.240 203.130 ;
        RECT 110.455 202.470 110.765 202.800 ;
        RECT 110.935 202.470 111.240 202.800 ;
        RECT 111.415 202.470 111.700 203.130 ;
        RECT 111.895 202.470 112.160 203.130 ;
        RECT 112.375 202.470 112.620 203.130 ;
        RECT 110.595 202.300 110.765 202.470 ;
        RECT 112.790 202.300 112.960 203.300 ;
        RECT 113.305 202.970 113.585 204.110 ;
        RECT 113.755 202.960 114.085 203.940 ;
        RECT 114.255 202.970 114.515 204.110 ;
        RECT 114.690 203.720 115.025 203.940 ;
        RECT 116.030 203.730 116.385 204.110 ;
        RECT 114.690 203.100 114.945 203.720 ;
        RECT 115.195 203.560 115.425 203.600 ;
        RECT 116.555 203.560 116.805 203.940 ;
        RECT 115.195 203.360 116.805 203.560 ;
        RECT 115.195 203.270 115.380 203.360 ;
        RECT 115.970 203.350 116.805 203.360 ;
        RECT 117.055 203.330 117.305 204.110 ;
        RECT 117.475 203.260 117.735 203.940 ;
        RECT 115.535 203.160 115.865 203.190 ;
        RECT 115.535 203.100 117.335 203.160 ;
        RECT 114.690 202.990 117.395 203.100 ;
        RECT 113.315 202.530 113.650 202.800 ;
        RECT 113.820 202.360 113.990 202.960 ;
        RECT 114.690 202.930 115.865 202.990 ;
        RECT 117.195 202.955 117.395 202.990 ;
        RECT 114.160 202.550 114.495 202.800 ;
        RECT 114.685 202.550 115.175 202.750 ;
        RECT 115.365 202.550 115.840 202.760 ;
        RECT 110.095 201.775 110.425 202.285 ;
        RECT 110.595 202.130 112.960 202.300 ;
        RECT 110.595 201.560 110.925 201.960 ;
        RECT 111.975 201.790 112.305 202.130 ;
        RECT 112.475 201.560 112.805 201.960 ;
        RECT 113.305 201.560 113.615 202.360 ;
        RECT 113.820 201.730 114.515 202.360 ;
        RECT 114.690 201.560 115.145 202.325 ;
        RECT 115.620 202.150 115.840 202.550 ;
        RECT 116.085 202.550 116.415 202.760 ;
        RECT 116.085 202.150 116.295 202.550 ;
        RECT 116.585 202.515 116.995 202.820 ;
        RECT 117.225 202.380 117.395 202.955 ;
        RECT 117.125 202.260 117.395 202.380 ;
        RECT 116.550 202.215 117.395 202.260 ;
        RECT 116.550 202.090 117.305 202.215 ;
        RECT 116.550 201.940 116.720 202.090 ;
        RECT 117.565 202.060 117.735 203.260 ;
        RECT 115.420 201.730 116.720 201.940 ;
        RECT 116.975 201.560 117.305 201.920 ;
        RECT 117.475 201.730 117.735 202.060 ;
        RECT 118.370 202.920 118.625 203.800 ;
        RECT 118.795 202.970 119.100 204.110 ;
        RECT 119.440 203.730 119.770 204.110 ;
        RECT 119.950 203.560 120.120 203.850 ;
        RECT 120.290 203.650 120.540 204.110 ;
        RECT 119.320 203.390 120.120 203.560 ;
        RECT 120.710 203.600 121.580 203.940 ;
        RECT 118.370 202.270 118.580 202.920 ;
        RECT 119.320 202.800 119.490 203.390 ;
        RECT 120.710 203.220 120.880 203.600 ;
        RECT 121.815 203.480 121.985 203.940 ;
        RECT 122.155 203.650 122.525 204.110 ;
        RECT 122.820 203.510 122.990 203.850 ;
        RECT 123.160 203.680 123.490 204.110 ;
        RECT 123.725 203.510 123.895 203.850 ;
        RECT 119.660 203.050 120.880 203.220 ;
        RECT 121.050 203.140 121.510 203.430 ;
        RECT 121.815 203.310 122.375 203.480 ;
        RECT 122.820 203.340 123.895 203.510 ;
        RECT 124.065 203.610 124.745 203.940 ;
        RECT 124.960 203.610 125.210 203.940 ;
        RECT 125.380 203.650 125.630 204.110 ;
        RECT 122.205 203.170 122.375 203.310 ;
        RECT 121.050 203.130 122.015 203.140 ;
        RECT 120.710 202.960 120.880 203.050 ;
        RECT 121.340 202.970 122.015 203.130 ;
        RECT 118.750 202.770 119.490 202.800 ;
        RECT 118.750 202.470 119.665 202.770 ;
        RECT 119.340 202.295 119.665 202.470 ;
        RECT 118.370 201.740 118.625 202.270 ;
        RECT 118.795 201.560 119.100 202.020 ;
        RECT 119.345 201.940 119.665 202.295 ;
        RECT 119.835 202.510 120.375 202.880 ;
        RECT 120.710 202.790 121.115 202.960 ;
        RECT 119.835 202.110 120.075 202.510 ;
        RECT 120.555 202.340 120.775 202.620 ;
        RECT 120.245 202.170 120.775 202.340 ;
        RECT 120.245 201.940 120.415 202.170 ;
        RECT 120.945 202.010 121.115 202.790 ;
        RECT 121.285 202.180 121.635 202.800 ;
        RECT 121.805 202.180 122.015 202.970 ;
        RECT 122.205 203.000 123.705 203.170 ;
        RECT 122.205 202.310 122.375 203.000 ;
        RECT 124.065 202.830 124.235 203.610 ;
        RECT 125.040 203.480 125.210 203.610 ;
        RECT 122.545 202.660 124.235 202.830 ;
        RECT 124.405 203.050 124.870 203.440 ;
        RECT 125.040 203.310 125.435 203.480 ;
        RECT 122.545 202.480 122.715 202.660 ;
        RECT 119.345 201.770 120.415 201.940 ;
        RECT 120.585 201.560 120.775 202.000 ;
        RECT 120.945 201.730 121.895 202.010 ;
        RECT 122.205 201.920 122.465 202.310 ;
        RECT 122.885 202.240 123.675 202.490 ;
        RECT 122.115 201.750 122.465 201.920 ;
        RECT 122.675 201.560 123.005 202.020 ;
        RECT 123.880 201.950 124.050 202.660 ;
        RECT 124.405 202.460 124.575 203.050 ;
        RECT 124.220 202.240 124.575 202.460 ;
        RECT 124.745 202.240 125.095 202.860 ;
        RECT 125.265 201.950 125.435 203.310 ;
        RECT 125.800 203.140 126.125 203.925 ;
        RECT 125.605 202.090 126.065 203.140 ;
        RECT 123.880 201.780 124.735 201.950 ;
        RECT 124.940 201.780 125.435 201.950 ;
        RECT 125.605 201.560 125.935 201.920 ;
        RECT 126.295 201.820 126.465 203.940 ;
        RECT 126.635 203.610 126.965 204.110 ;
        RECT 127.135 203.440 127.390 203.940 ;
        RECT 126.640 203.270 127.390 203.440 ;
        RECT 127.565 203.390 128.025 203.940 ;
        RECT 128.215 203.390 128.545 204.110 ;
        RECT 126.640 202.280 126.870 203.270 ;
        RECT 127.040 202.450 127.390 203.100 ;
        RECT 126.640 202.110 127.390 202.280 ;
        RECT 126.635 201.560 126.965 201.940 ;
        RECT 127.135 201.820 127.390 202.110 ;
        RECT 127.565 202.020 127.815 203.390 ;
        RECT 128.745 203.220 129.045 203.770 ;
        RECT 129.215 203.440 129.495 204.110 ;
        RECT 128.105 203.050 129.045 203.220 ;
        RECT 128.105 202.800 128.275 203.050 ;
        RECT 129.415 202.800 129.680 203.160 ;
        RECT 129.865 202.945 130.155 204.110 ;
        RECT 127.985 202.470 128.275 202.800 ;
        RECT 128.445 202.550 128.785 202.800 ;
        RECT 129.005 202.550 129.680 202.800 ;
        RECT 130.330 202.920 130.585 203.800 ;
        RECT 130.755 202.970 131.060 204.110 ;
        RECT 131.400 203.730 131.730 204.110 ;
        RECT 131.910 203.560 132.080 203.850 ;
        RECT 132.250 203.650 132.500 204.110 ;
        RECT 131.280 203.390 132.080 203.560 ;
        RECT 132.670 203.600 133.540 203.940 ;
        RECT 128.105 202.380 128.275 202.470 ;
        RECT 128.105 202.190 129.495 202.380 ;
        RECT 127.565 201.730 128.125 202.020 ;
        RECT 128.295 201.560 128.545 202.020 ;
        RECT 129.165 201.830 129.495 202.190 ;
        RECT 129.865 201.560 130.155 202.285 ;
        RECT 130.330 202.270 130.540 202.920 ;
        RECT 131.280 202.800 131.450 203.390 ;
        RECT 132.670 203.220 132.840 203.600 ;
        RECT 133.775 203.480 133.945 203.940 ;
        RECT 134.115 203.650 134.485 204.110 ;
        RECT 134.780 203.510 134.950 203.850 ;
        RECT 135.120 203.680 135.450 204.110 ;
        RECT 135.685 203.510 135.855 203.850 ;
        RECT 131.620 203.050 132.840 203.220 ;
        RECT 133.010 203.140 133.470 203.430 ;
        RECT 133.775 203.310 134.335 203.480 ;
        RECT 134.780 203.340 135.855 203.510 ;
        RECT 136.025 203.610 136.705 203.940 ;
        RECT 136.920 203.610 137.170 203.940 ;
        RECT 137.340 203.650 137.590 204.110 ;
        RECT 134.165 203.170 134.335 203.310 ;
        RECT 133.010 203.130 133.975 203.140 ;
        RECT 132.670 202.960 132.840 203.050 ;
        RECT 133.300 202.970 133.975 203.130 ;
        RECT 130.710 202.770 131.450 202.800 ;
        RECT 130.710 202.470 131.625 202.770 ;
        RECT 131.300 202.295 131.625 202.470 ;
        RECT 130.330 201.740 130.585 202.270 ;
        RECT 130.755 201.560 131.060 202.020 ;
        RECT 131.305 201.940 131.625 202.295 ;
        RECT 131.795 202.510 132.335 202.880 ;
        RECT 132.670 202.790 133.075 202.960 ;
        RECT 131.795 202.110 132.035 202.510 ;
        RECT 132.515 202.340 132.735 202.620 ;
        RECT 132.205 202.170 132.735 202.340 ;
        RECT 132.205 201.940 132.375 202.170 ;
        RECT 132.905 202.010 133.075 202.790 ;
        RECT 133.245 202.180 133.595 202.800 ;
        RECT 133.765 202.180 133.975 202.970 ;
        RECT 134.165 203.000 135.665 203.170 ;
        RECT 134.165 202.310 134.335 203.000 ;
        RECT 136.025 202.830 136.195 203.610 ;
        RECT 137.000 203.480 137.170 203.610 ;
        RECT 134.505 202.660 136.195 202.830 ;
        RECT 136.365 203.050 136.830 203.440 ;
        RECT 137.000 203.310 137.395 203.480 ;
        RECT 134.505 202.480 134.675 202.660 ;
        RECT 131.305 201.770 132.375 201.940 ;
        RECT 132.545 201.560 132.735 202.000 ;
        RECT 132.905 201.730 133.855 202.010 ;
        RECT 134.165 201.920 134.425 202.310 ;
        RECT 134.845 202.240 135.635 202.490 ;
        RECT 134.075 201.750 134.425 201.920 ;
        RECT 134.635 201.560 134.965 202.020 ;
        RECT 135.840 201.950 136.010 202.660 ;
        RECT 136.365 202.460 136.535 203.050 ;
        RECT 136.180 202.240 136.535 202.460 ;
        RECT 136.705 202.240 137.055 202.860 ;
        RECT 137.225 201.950 137.395 203.310 ;
        RECT 137.760 203.140 138.085 203.925 ;
        RECT 137.565 202.090 138.025 203.140 ;
        RECT 135.840 201.780 136.695 201.950 ;
        RECT 136.900 201.780 137.395 201.950 ;
        RECT 137.565 201.560 137.895 201.920 ;
        RECT 138.255 201.820 138.425 203.940 ;
        RECT 138.595 203.610 138.925 204.110 ;
        RECT 139.095 203.440 139.350 203.940 ;
        RECT 138.600 203.270 139.350 203.440 ;
        RECT 138.600 202.280 138.830 203.270 ;
        RECT 139.000 202.450 139.350 203.100 ;
        RECT 139.565 202.970 139.795 204.110 ;
        RECT 139.965 202.960 140.295 203.940 ;
        RECT 140.465 202.970 140.675 204.110 ;
        RECT 141.455 203.180 141.625 203.940 ;
        RECT 141.805 203.350 142.135 204.110 ;
        RECT 141.455 203.010 142.120 203.180 ;
        RECT 142.305 203.035 142.575 203.940 ;
        RECT 139.545 202.550 139.875 202.800 ;
        RECT 138.600 202.110 139.350 202.280 ;
        RECT 138.595 201.560 138.925 201.940 ;
        RECT 139.095 201.820 139.350 202.110 ;
        RECT 139.565 201.560 139.795 202.380 ;
        RECT 140.045 202.360 140.295 202.960 ;
        RECT 141.950 202.865 142.120 203.010 ;
        RECT 141.385 202.460 141.715 202.830 ;
        RECT 141.950 202.535 142.235 202.865 ;
        RECT 139.965 201.730 140.295 202.360 ;
        RECT 140.465 201.560 140.675 202.380 ;
        RECT 141.950 202.280 142.120 202.535 ;
        RECT 141.455 202.110 142.120 202.280 ;
        RECT 142.405 202.235 142.575 203.035 ;
        RECT 142.835 203.180 143.005 203.940 ;
        RECT 143.220 203.350 143.550 204.110 ;
        RECT 142.835 203.010 143.550 203.180 ;
        RECT 143.720 203.035 143.975 203.940 ;
        RECT 142.745 202.460 143.100 202.830 ;
        RECT 143.380 202.800 143.550 203.010 ;
        RECT 143.380 202.470 143.635 202.800 ;
        RECT 143.380 202.280 143.550 202.470 ;
        RECT 143.805 202.305 143.975 203.035 ;
        RECT 144.150 202.960 144.410 204.110 ;
        RECT 144.675 203.180 144.845 203.940 ;
        RECT 145.060 203.350 145.390 204.110 ;
        RECT 144.675 203.010 145.390 203.180 ;
        RECT 145.560 203.035 145.815 203.940 ;
        RECT 144.585 202.460 144.940 202.830 ;
        RECT 145.220 202.800 145.390 203.010 ;
        RECT 145.220 202.470 145.475 202.800 ;
        RECT 141.455 201.730 141.625 202.110 ;
        RECT 141.805 201.560 142.135 201.940 ;
        RECT 142.315 201.730 142.575 202.235 ;
        RECT 142.835 202.110 143.550 202.280 ;
        RECT 142.835 201.730 143.005 202.110 ;
        RECT 143.220 201.560 143.550 201.940 ;
        RECT 143.720 201.730 143.975 202.305 ;
        RECT 144.150 201.560 144.410 202.400 ;
        RECT 145.220 202.280 145.390 202.470 ;
        RECT 145.645 202.305 145.815 203.035 ;
        RECT 145.990 202.960 146.250 204.110 ;
        RECT 146.425 203.020 147.635 204.110 ;
        RECT 146.425 202.480 146.945 203.020 ;
        RECT 144.675 202.110 145.390 202.280 ;
        RECT 144.675 201.730 144.845 202.110 ;
        RECT 145.060 201.560 145.390 201.940 ;
        RECT 145.560 201.730 145.815 202.305 ;
        RECT 145.990 201.560 146.250 202.400 ;
        RECT 147.115 202.310 147.635 202.850 ;
        RECT 146.425 201.560 147.635 202.310 ;
        RECT 13.860 201.390 147.720 201.560 ;
        RECT 13.945 200.640 15.155 201.390 ;
        RECT 13.945 200.100 14.465 200.640 ;
        RECT 15.330 200.550 15.590 201.390 ;
        RECT 15.765 200.645 16.020 201.220 ;
        RECT 16.190 201.010 16.520 201.390 ;
        RECT 16.735 200.840 16.905 201.220 ;
        RECT 16.190 200.670 16.905 200.840 ;
        RECT 14.635 199.930 15.155 200.470 ;
        RECT 13.945 198.840 15.155 199.930 ;
        RECT 15.330 198.840 15.590 199.990 ;
        RECT 15.765 199.915 15.935 200.645 ;
        RECT 16.190 200.480 16.360 200.670 ;
        RECT 17.170 200.550 17.430 201.390 ;
        RECT 17.605 200.645 17.860 201.220 ;
        RECT 18.030 201.010 18.360 201.390 ;
        RECT 18.575 200.840 18.745 201.220 ;
        RECT 18.030 200.670 18.745 200.840 ;
        RECT 19.470 200.840 19.725 201.130 ;
        RECT 19.895 201.010 20.225 201.390 ;
        RECT 19.470 200.670 20.220 200.840 ;
        RECT 16.105 200.150 16.360 200.480 ;
        RECT 16.190 199.940 16.360 200.150 ;
        RECT 16.640 200.120 16.995 200.490 ;
        RECT 15.765 199.010 16.020 199.915 ;
        RECT 16.190 199.770 16.905 199.940 ;
        RECT 16.190 198.840 16.520 199.600 ;
        RECT 16.735 199.010 16.905 199.770 ;
        RECT 17.170 198.840 17.430 199.990 ;
        RECT 17.605 199.915 17.775 200.645 ;
        RECT 18.030 200.480 18.200 200.670 ;
        RECT 17.945 200.150 18.200 200.480 ;
        RECT 18.030 199.940 18.200 200.150 ;
        RECT 18.480 200.120 18.835 200.490 ;
        RECT 17.605 199.010 17.860 199.915 ;
        RECT 18.030 199.770 18.745 199.940 ;
        RECT 19.470 199.850 19.820 200.500 ;
        RECT 18.030 198.840 18.360 199.600 ;
        RECT 18.575 199.010 18.745 199.770 ;
        RECT 19.990 199.680 20.220 200.670 ;
        RECT 19.470 199.510 20.220 199.680 ;
        RECT 19.470 199.010 19.725 199.510 ;
        RECT 19.895 198.840 20.225 199.340 ;
        RECT 20.395 199.010 20.565 201.130 ;
        RECT 20.925 201.030 21.255 201.390 ;
        RECT 21.425 201.000 21.920 201.170 ;
        RECT 22.125 201.000 22.980 201.170 ;
        RECT 20.795 199.810 21.255 200.860 ;
        RECT 20.735 199.025 21.060 199.810 ;
        RECT 21.425 199.640 21.595 201.000 ;
        RECT 21.765 200.090 22.115 200.710 ;
        RECT 22.285 200.490 22.640 200.710 ;
        RECT 22.285 199.900 22.455 200.490 ;
        RECT 22.810 200.290 22.980 201.000 ;
        RECT 23.855 200.930 24.185 201.390 ;
        RECT 24.395 201.030 24.745 201.200 ;
        RECT 23.185 200.460 23.975 200.710 ;
        RECT 24.395 200.640 24.655 201.030 ;
        RECT 24.965 200.940 25.915 201.220 ;
        RECT 26.085 200.950 26.275 201.390 ;
        RECT 26.445 201.010 27.515 201.180 ;
        RECT 24.145 200.290 24.315 200.470 ;
        RECT 21.425 199.470 21.820 199.640 ;
        RECT 21.990 199.510 22.455 199.900 ;
        RECT 22.625 200.120 24.315 200.290 ;
        RECT 21.650 199.340 21.820 199.470 ;
        RECT 22.625 199.340 22.795 200.120 ;
        RECT 24.485 199.950 24.655 200.640 ;
        RECT 23.155 199.780 24.655 199.950 ;
        RECT 24.845 199.980 25.055 200.770 ;
        RECT 25.225 200.150 25.575 200.770 ;
        RECT 25.745 200.160 25.915 200.940 ;
        RECT 26.445 200.780 26.615 201.010 ;
        RECT 26.085 200.610 26.615 200.780 ;
        RECT 26.085 200.330 26.305 200.610 ;
        RECT 26.785 200.440 27.025 200.840 ;
        RECT 25.745 199.990 26.150 200.160 ;
        RECT 26.485 200.070 27.025 200.440 ;
        RECT 27.195 200.655 27.515 201.010 ;
        RECT 27.195 200.400 27.520 200.655 ;
        RECT 27.715 200.580 27.885 201.390 ;
        RECT 28.055 200.740 28.385 201.220 ;
        RECT 28.555 200.920 28.725 201.390 ;
        RECT 28.895 200.740 29.225 201.220 ;
        RECT 29.395 200.920 29.565 201.390 ;
        RECT 30.705 200.760 31.035 201.120 ;
        RECT 31.655 200.930 31.905 201.390 ;
        RECT 32.075 200.930 32.635 201.220 ;
        RECT 28.055 200.570 29.820 200.740 ;
        RECT 30.705 200.570 32.095 200.760 ;
        RECT 27.195 200.190 29.225 200.400 ;
        RECT 27.195 200.180 27.540 200.190 ;
        RECT 24.845 199.820 25.520 199.980 ;
        RECT 25.980 199.900 26.150 199.990 ;
        RECT 24.845 199.810 25.810 199.820 ;
        RECT 24.485 199.640 24.655 199.780 ;
        RECT 21.230 198.840 21.480 199.300 ;
        RECT 21.650 199.010 21.900 199.340 ;
        RECT 22.115 199.010 22.795 199.340 ;
        RECT 22.965 199.440 24.040 199.610 ;
        RECT 24.485 199.470 25.045 199.640 ;
        RECT 25.350 199.520 25.810 199.810 ;
        RECT 25.980 199.730 27.200 199.900 ;
        RECT 22.965 199.100 23.135 199.440 ;
        RECT 23.370 198.840 23.700 199.270 ;
        RECT 23.870 199.100 24.040 199.440 ;
        RECT 24.335 198.840 24.705 199.300 ;
        RECT 24.875 199.010 25.045 199.470 ;
        RECT 25.980 199.350 26.150 199.730 ;
        RECT 27.370 199.560 27.540 200.180 ;
        RECT 29.410 200.020 29.820 200.570 ;
        RECT 31.925 200.480 32.095 200.570 ;
        RECT 25.280 199.010 26.150 199.350 ;
        RECT 26.740 199.390 27.540 199.560 ;
        RECT 26.320 198.840 26.570 199.300 ;
        RECT 26.740 199.100 26.910 199.390 ;
        RECT 27.090 198.840 27.420 199.220 ;
        RECT 27.715 198.840 27.885 199.900 ;
        RECT 28.095 199.850 29.820 200.020 ;
        RECT 30.520 200.150 31.195 200.400 ;
        RECT 31.415 200.150 31.755 200.400 ;
        RECT 31.925 200.150 32.215 200.480 ;
        RECT 28.095 199.010 28.385 199.850 ;
        RECT 28.555 198.840 28.725 199.680 ;
        RECT 28.935 199.010 29.185 199.850 ;
        RECT 30.520 199.790 30.785 200.150 ;
        RECT 31.925 199.900 32.095 200.150 ;
        RECT 31.155 199.730 32.095 199.900 ;
        RECT 29.395 198.840 29.565 199.680 ;
        RECT 30.705 198.840 30.985 199.510 ;
        RECT 31.155 199.180 31.455 199.730 ;
        RECT 32.385 199.560 32.635 200.930 ;
        RECT 32.970 200.880 33.210 201.390 ;
        RECT 33.390 200.880 33.670 201.210 ;
        RECT 33.900 200.880 34.115 201.390 ;
        RECT 32.865 200.150 33.220 200.710 ;
        RECT 33.390 199.980 33.560 200.880 ;
        RECT 33.730 200.150 33.995 200.710 ;
        RECT 34.285 200.650 34.900 201.220 ;
        RECT 34.245 199.980 34.415 200.480 ;
        RECT 32.990 199.810 34.415 199.980 ;
        RECT 32.990 199.635 33.380 199.810 ;
        RECT 31.655 198.840 31.985 199.560 ;
        RECT 32.175 199.010 32.635 199.560 ;
        RECT 33.865 198.840 34.195 199.640 ;
        RECT 34.585 199.630 34.900 200.650 ;
        RECT 34.365 199.010 34.900 199.630 ;
        RECT 35.125 200.890 35.380 201.220 ;
        RECT 35.595 200.910 35.925 201.390 ;
        RECT 36.095 200.970 37.630 201.220 ;
        RECT 35.125 200.810 35.310 200.890 ;
        RECT 35.125 199.680 35.295 200.810 ;
        RECT 36.095 200.740 36.265 200.970 ;
        RECT 35.465 200.570 36.265 200.740 ;
        RECT 35.465 200.020 35.635 200.570 ;
        RECT 36.445 200.400 36.730 200.800 ;
        RECT 35.865 200.370 36.230 200.400 ;
        RECT 35.855 200.200 36.230 200.370 ;
        RECT 36.400 200.200 36.730 200.400 ;
        RECT 37.000 200.400 37.280 200.800 ;
        RECT 37.460 200.740 37.630 200.970 ;
        RECT 37.855 200.910 38.185 201.390 ;
        RECT 38.355 200.740 38.525 201.220 ;
        RECT 37.460 200.570 38.525 200.740 ;
        RECT 39.705 200.665 39.995 201.390 ;
        RECT 40.185 200.890 40.440 201.220 ;
        RECT 40.655 200.910 40.985 201.390 ;
        RECT 41.155 200.970 42.690 201.220 ;
        RECT 40.185 200.880 40.395 200.890 ;
        RECT 40.185 200.810 40.370 200.880 ;
        RECT 37.000 200.200 37.475 200.400 ;
        RECT 37.645 200.200 38.090 200.400 ;
        RECT 38.260 200.190 38.610 200.400 ;
        RECT 35.465 199.850 38.525 200.020 ;
        RECT 35.125 199.010 35.380 199.680 ;
        RECT 35.550 198.840 35.880 199.600 ;
        RECT 36.050 199.440 37.685 199.680 ;
        RECT 36.050 199.010 36.300 199.440 ;
        RECT 37.455 199.350 37.685 199.440 ;
        RECT 36.470 198.840 36.825 199.260 ;
        RECT 37.015 199.180 37.345 199.220 ;
        RECT 37.855 199.180 38.185 199.680 ;
        RECT 37.015 199.010 38.185 199.180 ;
        RECT 38.355 199.010 38.525 199.850 ;
        RECT 39.705 198.840 39.995 200.005 ;
        RECT 40.185 199.680 40.355 200.810 ;
        RECT 41.155 200.740 41.325 200.970 ;
        RECT 40.525 200.570 41.325 200.740 ;
        RECT 40.525 200.020 40.695 200.570 ;
        RECT 41.505 200.400 41.790 200.800 ;
        RECT 40.925 200.200 41.290 200.400 ;
        RECT 41.460 200.200 41.790 200.400 ;
        RECT 42.060 200.400 42.340 200.800 ;
        RECT 42.520 200.740 42.690 200.970 ;
        RECT 42.915 200.910 43.245 201.390 ;
        RECT 43.415 200.740 43.585 201.220 ;
        RECT 42.520 200.570 43.585 200.740 ;
        RECT 43.880 200.650 44.495 201.220 ;
        RECT 44.665 200.880 44.880 201.390 ;
        RECT 45.110 200.880 45.390 201.210 ;
        RECT 45.570 200.880 45.810 201.390 ;
        RECT 42.060 200.200 42.535 200.400 ;
        RECT 42.705 200.200 43.150 200.400 ;
        RECT 43.320 200.190 43.670 200.400 ;
        RECT 40.525 199.850 43.585 200.020 ;
        RECT 40.185 199.010 40.440 199.680 ;
        RECT 40.610 198.840 40.940 199.600 ;
        RECT 41.110 199.440 42.745 199.680 ;
        RECT 41.110 199.010 41.360 199.440 ;
        RECT 42.515 199.350 42.745 199.440 ;
        RECT 41.530 198.840 41.885 199.260 ;
        RECT 42.075 199.180 42.405 199.220 ;
        RECT 42.915 199.180 43.245 199.680 ;
        RECT 42.075 199.010 43.245 199.180 ;
        RECT 43.415 199.010 43.585 199.850 ;
        RECT 43.880 199.630 44.195 200.650 ;
        RECT 44.365 199.980 44.535 200.480 ;
        RECT 44.785 200.150 45.050 200.710 ;
        RECT 45.220 199.980 45.390 200.880 ;
        RECT 45.560 200.150 45.915 200.710 ;
        RECT 46.165 200.580 46.405 201.390 ;
        RECT 46.575 200.580 46.905 201.220 ;
        RECT 47.075 200.580 47.345 201.390 ;
        RECT 46.145 200.150 46.495 200.400 ;
        RECT 46.665 199.980 46.835 200.580 ;
        RECT 47.005 200.150 47.355 200.400 ;
        RECT 44.365 199.810 45.790 199.980 ;
        RECT 43.880 199.010 44.415 199.630 ;
        RECT 44.585 198.840 44.915 199.640 ;
        RECT 45.400 199.635 45.790 199.810 ;
        RECT 46.155 199.810 46.835 199.980 ;
        RECT 46.155 199.025 46.485 199.810 ;
        RECT 47.015 198.840 47.345 199.980 ;
        RECT 47.530 199.790 47.865 201.210 ;
        RECT 48.045 201.020 48.790 201.390 ;
        RECT 49.355 200.850 49.610 201.210 ;
        RECT 49.790 201.020 50.120 201.390 ;
        RECT 50.300 200.850 50.525 201.210 ;
        RECT 48.040 200.660 50.525 200.850 ;
        RECT 48.040 199.970 48.265 200.660 ;
        RECT 50.785 200.570 51.015 201.390 ;
        RECT 51.185 200.590 51.515 201.220 ;
        RECT 48.465 200.150 48.745 200.480 ;
        RECT 48.925 200.150 49.500 200.480 ;
        RECT 49.680 200.150 50.115 200.480 ;
        RECT 50.295 200.150 50.565 200.480 ;
        RECT 50.765 200.150 51.095 200.400 ;
        RECT 51.265 199.990 51.515 200.590 ;
        RECT 51.685 200.570 51.895 201.390 ;
        RECT 52.165 200.570 52.395 201.390 ;
        RECT 52.565 200.590 52.895 201.220 ;
        RECT 52.145 200.150 52.475 200.400 ;
        RECT 52.645 199.990 52.895 200.590 ;
        RECT 53.065 200.570 53.275 201.390 ;
        RECT 54.435 200.580 54.705 201.390 ;
        RECT 54.875 200.580 55.205 201.220 ;
        RECT 55.375 200.580 55.615 201.390 ;
        RECT 55.970 200.880 56.210 201.390 ;
        RECT 56.390 200.880 56.670 201.210 ;
        RECT 56.900 200.880 57.115 201.390 ;
        RECT 54.425 200.150 54.775 200.400 ;
        RECT 48.040 199.790 50.535 199.970 ;
        RECT 47.530 199.020 47.795 199.790 ;
        RECT 47.965 198.840 48.295 199.560 ;
        RECT 48.485 199.380 49.675 199.610 ;
        RECT 48.485 199.020 48.745 199.380 ;
        RECT 48.915 198.840 49.245 199.210 ;
        RECT 49.415 199.020 49.675 199.380 ;
        RECT 50.245 199.020 50.535 199.790 ;
        RECT 50.785 198.840 51.015 199.980 ;
        RECT 51.185 199.010 51.515 199.990 ;
        RECT 51.685 198.840 51.895 199.980 ;
        RECT 52.165 198.840 52.395 199.980 ;
        RECT 52.565 199.010 52.895 199.990 ;
        RECT 54.945 199.980 55.115 200.580 ;
        RECT 55.285 200.150 55.635 200.400 ;
        RECT 55.865 200.150 56.220 200.710 ;
        RECT 56.390 199.980 56.560 200.880 ;
        RECT 56.730 200.150 56.995 200.710 ;
        RECT 57.285 200.650 57.900 201.220 ;
        RECT 57.245 199.980 57.415 200.480 ;
        RECT 53.065 198.840 53.275 199.980 ;
        RECT 54.435 198.840 54.765 199.980 ;
        RECT 54.945 199.810 55.625 199.980 ;
        RECT 55.295 199.025 55.625 199.810 ;
        RECT 55.990 199.810 57.415 199.980 ;
        RECT 55.990 199.635 56.380 199.810 ;
        RECT 56.865 198.840 57.195 199.640 ;
        RECT 57.585 199.630 57.900 200.650 ;
        RECT 58.195 200.740 58.365 201.220 ;
        RECT 58.535 200.910 58.865 201.390 ;
        RECT 59.090 200.970 60.625 201.220 ;
        RECT 59.090 200.740 59.260 200.970 ;
        RECT 58.195 200.570 59.260 200.740 ;
        RECT 59.440 200.400 59.720 200.800 ;
        RECT 58.110 200.190 58.460 200.400 ;
        RECT 58.630 200.200 59.075 200.400 ;
        RECT 59.245 200.200 59.720 200.400 ;
        RECT 59.990 200.400 60.275 200.800 ;
        RECT 60.455 200.740 60.625 200.970 ;
        RECT 60.795 200.910 61.125 201.390 ;
        RECT 61.340 200.890 61.595 201.220 ;
        RECT 61.410 200.810 61.595 200.890 ;
        RECT 60.455 200.570 61.255 200.740 ;
        RECT 59.990 200.200 60.320 200.400 ;
        RECT 60.490 200.370 60.855 200.400 ;
        RECT 60.490 200.200 60.865 200.370 ;
        RECT 61.085 200.020 61.255 200.570 ;
        RECT 57.365 199.010 57.900 199.630 ;
        RECT 58.195 199.850 61.255 200.020 ;
        RECT 58.195 199.010 58.365 199.850 ;
        RECT 61.425 199.690 61.595 200.810 ;
        RECT 61.385 199.680 61.595 199.690 ;
        RECT 58.535 199.180 58.865 199.680 ;
        RECT 59.035 199.440 60.670 199.680 ;
        RECT 59.035 199.350 59.265 199.440 ;
        RECT 59.375 199.180 59.705 199.220 ;
        RECT 58.535 199.010 59.705 199.180 ;
        RECT 59.895 198.840 60.250 199.260 ;
        RECT 60.420 199.010 60.670 199.440 ;
        RECT 60.840 198.840 61.170 199.600 ;
        RECT 61.340 199.010 61.595 199.680 ;
        RECT 61.795 199.020 62.055 201.210 ;
        RECT 62.315 201.020 62.985 201.390 ;
        RECT 63.165 200.840 63.475 201.210 ;
        RECT 62.245 200.640 63.475 200.840 ;
        RECT 62.245 199.970 62.535 200.640 ;
        RECT 63.655 200.460 63.885 201.100 ;
        RECT 64.065 200.660 64.355 201.390 ;
        RECT 65.465 200.665 65.755 201.390 ;
        RECT 62.715 200.150 63.180 200.460 ;
        RECT 63.360 200.150 63.885 200.460 ;
        RECT 64.065 200.150 64.365 200.480 ;
        RECT 62.245 199.750 63.015 199.970 ;
        RECT 62.225 198.840 62.565 199.570 ;
        RECT 62.745 199.020 63.015 199.750 ;
        RECT 63.195 199.730 64.355 199.970 ;
        RECT 63.195 199.020 63.425 199.730 ;
        RECT 63.595 198.840 63.925 199.550 ;
        RECT 64.095 199.020 64.355 199.730 ;
        RECT 65.465 198.840 65.755 200.005 ;
        RECT 65.935 199.020 66.195 201.210 ;
        RECT 66.455 201.020 67.125 201.390 ;
        RECT 67.305 200.840 67.615 201.210 ;
        RECT 66.385 200.640 67.615 200.840 ;
        RECT 66.385 199.970 66.675 200.640 ;
        RECT 67.795 200.460 68.025 201.100 ;
        RECT 68.205 200.660 68.495 201.390 ;
        RECT 68.685 200.990 69.275 201.220 ;
        RECT 70.320 200.990 70.650 201.390 ;
        RECT 66.855 200.150 67.320 200.460 ;
        RECT 67.500 200.150 68.025 200.460 ;
        RECT 68.205 200.150 68.505 200.480 ;
        RECT 68.685 199.980 68.975 200.990 ;
        RECT 70.850 200.820 71.275 201.030 ;
        RECT 69.145 200.650 71.275 200.820 ;
        RECT 71.460 200.820 71.715 201.170 ;
        RECT 71.885 200.990 72.215 201.390 ;
        RECT 72.385 200.820 72.555 201.170 ;
        RECT 72.725 200.990 73.105 201.390 ;
        RECT 71.460 200.650 73.125 200.820 ;
        RECT 73.295 200.715 73.570 201.060 ;
        RECT 69.145 200.150 69.315 200.650 ;
        RECT 69.605 200.150 69.935 200.480 ;
        RECT 70.125 200.150 70.395 200.480 ;
        RECT 70.585 200.150 70.935 200.480 ;
        RECT 66.385 199.750 67.155 199.970 ;
        RECT 66.365 198.840 66.705 199.570 ;
        RECT 66.885 199.020 67.155 199.750 ;
        RECT 67.335 199.730 68.495 199.970 ;
        RECT 67.335 199.020 67.565 199.730 ;
        RECT 67.735 198.840 68.065 199.550 ;
        RECT 68.235 199.020 68.495 199.730 ;
        RECT 68.685 199.810 70.230 199.980 ;
        RECT 68.685 199.010 69.275 199.810 ;
        RECT 69.445 198.840 69.730 199.640 ;
        RECT 69.900 199.010 70.230 199.810 ;
        RECT 70.400 198.840 70.650 199.980 ;
        RECT 71.105 199.880 71.275 200.650 ;
        RECT 72.955 200.480 73.125 200.650 ;
        RECT 71.445 200.150 71.790 200.480 ;
        RECT 71.960 200.150 72.785 200.480 ;
        RECT 72.955 200.150 73.230 200.480 ;
        RECT 70.850 199.550 71.275 199.880 ;
        RECT 71.465 199.690 71.790 199.980 ;
        RECT 71.960 199.860 72.155 200.150 ;
        RECT 72.955 199.980 73.125 200.150 ;
        RECT 73.400 199.980 73.570 200.715 ;
        RECT 72.465 199.810 73.125 199.980 ;
        RECT 72.465 199.690 72.635 199.810 ;
        RECT 71.465 199.520 72.635 199.690 ;
        RECT 71.445 199.060 72.635 199.350 ;
        RECT 72.805 198.840 73.085 199.640 ;
        RECT 73.295 199.010 73.570 199.980 ;
        RECT 74.670 199.790 75.005 201.210 ;
        RECT 75.185 201.020 75.930 201.390 ;
        RECT 76.495 200.850 76.750 201.210 ;
        RECT 76.930 201.020 77.260 201.390 ;
        RECT 77.440 200.850 77.665 201.210 ;
        RECT 75.180 200.660 77.665 200.850 ;
        RECT 77.895 200.665 78.225 201.175 ;
        RECT 78.395 200.990 78.725 201.390 ;
        RECT 79.775 200.820 80.105 201.160 ;
        RECT 80.275 200.990 80.605 201.390 ;
        RECT 75.180 199.970 75.405 200.660 ;
        RECT 75.605 200.150 75.885 200.480 ;
        RECT 76.065 200.150 76.640 200.480 ;
        RECT 76.820 200.150 77.255 200.480 ;
        RECT 77.435 200.150 77.705 200.480 ;
        RECT 77.895 200.030 78.085 200.665 ;
        RECT 78.395 200.650 80.760 200.820 ;
        RECT 78.395 200.480 78.565 200.650 ;
        RECT 78.255 200.150 78.565 200.480 ;
        RECT 78.735 200.150 79.040 200.480 ;
        RECT 75.180 199.790 77.675 199.970 ;
        RECT 74.670 199.020 74.935 199.790 ;
        RECT 75.105 198.840 75.435 199.560 ;
        RECT 75.625 199.380 76.815 199.610 ;
        RECT 75.625 199.020 75.885 199.380 ;
        RECT 76.055 198.840 76.385 199.210 ;
        RECT 76.555 199.020 76.815 199.380 ;
        RECT 77.385 199.020 77.675 199.790 ;
        RECT 77.895 199.900 78.115 200.030 ;
        RECT 77.895 199.050 78.225 199.900 ;
        RECT 78.395 198.840 78.645 199.980 ;
        RECT 78.825 199.820 79.040 200.150 ;
        RECT 79.215 199.820 79.500 200.480 ;
        RECT 79.695 199.820 79.960 200.480 ;
        RECT 80.175 199.820 80.420 200.480 ;
        RECT 80.590 199.650 80.760 200.650 ;
        RECT 78.835 199.480 80.125 199.650 ;
        RECT 78.835 199.060 79.085 199.480 ;
        RECT 79.315 198.840 79.645 199.310 ;
        RECT 79.875 199.060 80.125 199.480 ;
        RECT 80.305 199.480 80.760 199.650 ;
        RECT 81.565 200.650 82.075 201.220 ;
        RECT 82.245 200.830 82.415 201.390 ;
        RECT 82.620 200.820 82.950 201.220 ;
        RECT 83.125 200.990 83.455 201.390 ;
        RECT 83.690 201.010 85.075 201.220 ;
        RECT 83.690 200.820 84.020 201.010 ;
        RECT 82.620 200.650 84.020 200.820 ;
        RECT 84.190 200.650 84.615 200.840 ;
        RECT 84.785 200.740 85.075 201.010 ;
        RECT 81.565 200.030 81.740 200.650 ;
        RECT 81.925 200.400 82.115 200.480 ;
        RECT 82.485 200.400 82.655 200.480 ;
        RECT 81.925 200.150 82.290 200.400 ;
        RECT 82.485 200.150 82.735 200.400 ;
        RECT 82.945 200.150 83.290 200.480 ;
        RECT 81.565 199.980 81.795 200.030 ;
        RECT 82.120 199.980 82.290 200.150 ;
        RECT 80.305 199.050 80.635 199.480 ;
        RECT 81.565 199.020 81.950 199.980 ;
        RECT 82.120 199.810 82.795 199.980 ;
        RECT 82.165 198.840 82.455 199.640 ;
        RECT 82.625 199.180 82.795 199.810 ;
        RECT 82.965 199.350 83.290 200.150 ;
        RECT 83.460 199.815 83.735 200.480 ;
        RECT 83.920 199.815 84.275 200.480 ;
        RECT 84.445 199.640 84.615 200.650 ;
        RECT 85.335 200.570 85.505 201.390 ;
        RECT 85.675 200.740 86.005 201.220 ;
        RECT 86.175 200.910 86.345 201.390 ;
        RECT 86.530 200.740 86.860 201.220 ;
        RECT 85.675 200.570 86.860 200.740 ;
        RECT 87.105 200.650 87.835 201.215 ;
        RECT 88.050 200.930 88.800 201.220 ;
        RECT 89.310 200.930 89.640 201.390 ;
        RECT 84.800 200.150 85.075 200.480 ;
        RECT 85.250 200.150 85.600 200.400 ;
        RECT 83.660 199.390 84.615 199.640 ;
        RECT 83.660 199.180 83.990 199.390 ;
        RECT 82.625 199.010 83.990 199.180 ;
        RECT 84.785 198.840 85.075 199.980 ;
        RECT 85.250 198.840 85.600 199.980 ;
        RECT 85.770 199.010 86.215 200.400 ;
        RECT 86.385 200.150 86.860 200.400 ;
        RECT 86.620 199.070 86.860 200.150 ;
        RECT 87.105 199.010 87.320 200.650 ;
        RECT 87.490 200.150 87.835 200.480 ;
        RECT 87.490 198.840 87.835 199.980 ;
        RECT 88.050 199.640 88.420 200.930 ;
        RECT 89.860 200.740 90.130 200.950 ;
        RECT 88.795 200.570 90.130 200.740 ;
        RECT 91.225 200.665 91.515 201.390 ;
        RECT 91.685 200.650 92.125 201.220 ;
        RECT 92.295 200.880 93.665 201.050 ;
        RECT 93.835 200.990 94.165 201.390 ;
        RECT 88.795 200.400 88.965 200.570 ;
        RECT 88.590 200.150 88.965 200.400 ;
        RECT 89.135 200.160 89.610 200.400 ;
        RECT 89.780 200.160 90.130 200.400 ;
        RECT 88.795 199.980 88.965 200.150 ;
        RECT 91.685 200.030 91.895 200.650 ;
        RECT 92.295 200.480 92.465 200.880 ;
        RECT 93.485 200.820 93.665 200.880 ;
        RECT 94.345 200.820 94.735 201.030 ;
        RECT 92.065 200.150 92.465 200.480 ;
        RECT 92.635 200.150 92.895 200.710 ;
        RECT 93.065 200.150 93.315 200.710 ;
        RECT 93.485 200.650 94.735 200.820 ;
        RECT 93.585 200.150 93.855 200.480 ;
        RECT 94.045 200.150 94.395 200.480 ;
        RECT 88.795 199.810 90.130 199.980 ;
        RECT 89.850 199.650 90.130 199.810 ;
        RECT 88.050 199.470 89.220 199.640 ;
        RECT 88.505 198.840 88.720 199.300 ;
        RECT 88.890 199.010 89.220 199.470 ;
        RECT 89.390 198.840 89.640 199.640 ;
        RECT 91.225 198.840 91.515 200.005 ;
        RECT 91.685 199.980 91.915 200.030 ;
        RECT 91.685 199.810 93.690 199.980 ;
        RECT 91.900 198.840 92.115 199.640 ;
        RECT 92.405 199.010 92.735 199.810 ;
        RECT 92.905 198.840 93.190 199.640 ;
        RECT 93.360 199.010 93.690 199.810 ;
        RECT 93.860 198.840 94.110 199.980 ;
        RECT 94.565 199.880 94.735 200.650 ;
        RECT 94.905 200.620 96.575 201.390 ;
        RECT 97.210 200.625 97.665 201.390 ;
        RECT 97.940 201.010 99.240 201.220 ;
        RECT 99.495 201.030 99.825 201.390 ;
        RECT 99.070 200.860 99.240 201.010 ;
        RECT 99.995 200.890 100.255 201.220 ;
        RECT 94.905 200.100 95.655 200.620 ;
        RECT 95.825 199.930 96.575 200.450 ;
        RECT 98.140 200.400 98.360 200.800 ;
        RECT 97.205 200.200 97.695 200.400 ;
        RECT 97.885 200.190 98.360 200.400 ;
        RECT 98.605 200.400 98.815 200.800 ;
        RECT 99.070 200.735 99.825 200.860 ;
        RECT 99.070 200.690 99.915 200.735 ;
        RECT 99.645 200.570 99.915 200.690 ;
        RECT 98.605 200.190 98.935 200.400 ;
        RECT 99.105 200.130 99.515 200.435 ;
        RECT 94.310 199.550 94.735 199.880 ;
        RECT 94.905 198.840 96.575 199.930 ;
        RECT 97.210 199.960 98.385 200.020 ;
        RECT 99.745 199.995 99.915 200.570 ;
        RECT 99.715 199.960 99.915 199.995 ;
        RECT 97.210 199.850 99.915 199.960 ;
        RECT 97.210 199.230 97.465 199.850 ;
        RECT 98.055 199.790 99.855 199.850 ;
        RECT 98.055 199.760 98.385 199.790 ;
        RECT 100.085 199.690 100.255 200.890 ;
        RECT 100.425 200.640 101.635 201.390 ;
        RECT 100.425 200.100 100.945 200.640 ;
        RECT 101.805 200.590 102.500 201.220 ;
        RECT 102.705 200.590 103.015 201.390 ;
        RECT 103.185 200.590 103.880 201.220 ;
        RECT 104.085 200.590 104.395 201.390 ;
        RECT 104.570 200.625 105.025 201.390 ;
        RECT 105.300 201.010 106.600 201.220 ;
        RECT 106.855 201.030 107.185 201.390 ;
        RECT 106.430 200.860 106.600 201.010 ;
        RECT 107.355 200.890 107.615 201.220 ;
        RECT 101.115 199.930 101.635 200.470 ;
        RECT 101.825 200.150 102.160 200.400 ;
        RECT 102.330 200.030 102.500 200.590 ;
        RECT 102.670 200.150 103.005 200.420 ;
        RECT 103.205 200.150 103.540 200.400 ;
        RECT 102.325 199.990 102.500 200.030 ;
        RECT 103.710 199.990 103.880 200.590 ;
        RECT 104.050 200.150 104.385 200.420 ;
        RECT 105.500 200.400 105.720 200.800 ;
        RECT 104.565 200.200 105.055 200.400 ;
        RECT 105.245 200.190 105.720 200.400 ;
        RECT 105.965 200.400 106.175 200.800 ;
        RECT 106.430 200.735 107.185 200.860 ;
        RECT 106.430 200.690 107.275 200.735 ;
        RECT 107.005 200.570 107.275 200.690 ;
        RECT 105.965 200.190 106.295 200.400 ;
        RECT 106.465 200.130 106.875 200.435 ;
        RECT 97.715 199.590 97.900 199.680 ;
        RECT 98.490 199.590 99.325 199.600 ;
        RECT 97.715 199.390 99.325 199.590 ;
        RECT 97.715 199.350 97.945 199.390 ;
        RECT 97.210 199.010 97.545 199.230 ;
        RECT 98.550 198.840 98.905 199.220 ;
        RECT 99.075 199.010 99.325 199.390 ;
        RECT 99.575 198.840 99.825 199.620 ;
        RECT 99.995 199.010 100.255 199.690 ;
        RECT 100.425 198.840 101.635 199.930 ;
        RECT 101.805 198.840 102.065 199.980 ;
        RECT 102.235 199.010 102.565 199.990 ;
        RECT 102.735 198.840 103.015 199.980 ;
        RECT 103.185 198.840 103.445 199.980 ;
        RECT 103.615 199.010 103.945 199.990 ;
        RECT 104.115 198.840 104.395 199.980 ;
        RECT 104.570 199.960 105.745 200.020 ;
        RECT 107.105 199.995 107.275 200.570 ;
        RECT 107.075 199.960 107.275 199.995 ;
        RECT 104.570 199.850 107.275 199.960 ;
        RECT 104.570 199.230 104.825 199.850 ;
        RECT 105.415 199.790 107.215 199.850 ;
        RECT 105.415 199.760 105.745 199.790 ;
        RECT 107.445 199.690 107.615 200.890 ;
        RECT 107.785 200.880 108.090 201.390 ;
        RECT 107.785 200.150 108.100 200.710 ;
        RECT 108.270 200.400 108.520 201.210 ;
        RECT 108.690 200.865 108.950 201.390 ;
        RECT 109.130 200.400 109.380 201.210 ;
        RECT 109.550 200.830 109.810 201.390 ;
        RECT 109.980 200.740 110.240 201.195 ;
        RECT 110.410 200.910 110.670 201.390 ;
        RECT 110.840 200.740 111.100 201.195 ;
        RECT 111.270 200.910 111.530 201.390 ;
        RECT 111.700 200.740 111.960 201.195 ;
        RECT 112.130 200.910 112.375 201.390 ;
        RECT 112.545 200.740 112.820 201.195 ;
        RECT 112.990 200.910 113.235 201.390 ;
        RECT 113.405 200.740 113.665 201.195 ;
        RECT 113.845 200.910 114.095 201.390 ;
        RECT 114.265 200.740 114.525 201.195 ;
        RECT 114.705 200.910 114.955 201.390 ;
        RECT 115.125 200.740 115.385 201.195 ;
        RECT 115.565 200.910 115.825 201.390 ;
        RECT 115.995 200.740 116.255 201.195 ;
        RECT 116.425 200.910 116.725 201.390 ;
        RECT 109.980 200.570 116.725 200.740 ;
        RECT 116.985 200.665 117.275 201.390 ;
        RECT 118.480 200.760 118.765 201.220 ;
        RECT 118.935 200.930 119.205 201.390 ;
        RECT 118.480 200.590 119.435 200.760 ;
        RECT 108.270 200.150 115.390 200.400 ;
        RECT 105.075 199.590 105.260 199.680 ;
        RECT 105.850 199.590 106.685 199.600 ;
        RECT 105.075 199.390 106.685 199.590 ;
        RECT 105.075 199.350 105.305 199.390 ;
        RECT 104.570 199.010 104.905 199.230 ;
        RECT 105.910 198.840 106.265 199.220 ;
        RECT 106.435 199.010 106.685 199.390 ;
        RECT 106.935 198.840 107.185 199.620 ;
        RECT 107.355 199.010 107.615 199.690 ;
        RECT 107.795 198.840 108.090 199.650 ;
        RECT 108.270 199.010 108.515 200.150 ;
        RECT 108.690 198.840 108.950 199.650 ;
        RECT 109.130 199.015 109.380 200.150 ;
        RECT 115.560 199.980 116.725 200.570 ;
        RECT 109.980 199.755 116.725 199.980 ;
        RECT 109.980 199.740 115.385 199.755 ;
        RECT 109.550 198.845 109.810 199.640 ;
        RECT 109.980 199.015 110.240 199.740 ;
        RECT 110.410 198.845 110.670 199.570 ;
        RECT 110.840 199.015 111.100 199.740 ;
        RECT 111.270 198.845 111.530 199.570 ;
        RECT 111.700 199.015 111.960 199.740 ;
        RECT 112.130 198.845 112.390 199.570 ;
        RECT 112.560 199.015 112.820 199.740 ;
        RECT 112.990 198.845 113.235 199.570 ;
        RECT 113.405 199.015 113.665 199.740 ;
        RECT 113.850 198.845 114.095 199.570 ;
        RECT 114.265 199.015 114.525 199.740 ;
        RECT 114.710 198.845 114.955 199.570 ;
        RECT 115.125 199.015 115.385 199.740 ;
        RECT 115.570 198.845 115.825 199.570 ;
        RECT 115.995 199.015 116.285 199.755 ;
        RECT 109.550 198.840 115.825 198.845 ;
        RECT 116.455 198.840 116.725 199.585 ;
        RECT 116.985 198.840 117.275 200.005 ;
        RECT 118.365 199.860 119.055 200.420 ;
        RECT 119.225 199.690 119.435 200.590 ;
        RECT 118.480 199.470 119.435 199.690 ;
        RECT 119.605 200.420 120.005 201.220 ;
        RECT 120.195 200.760 120.475 201.220 ;
        RECT 120.995 200.930 121.320 201.390 ;
        RECT 120.195 200.590 121.320 200.760 ;
        RECT 121.490 200.650 121.875 201.220 ;
        RECT 120.870 200.480 121.320 200.590 ;
        RECT 119.605 199.860 120.700 200.420 ;
        RECT 120.870 200.150 121.425 200.480 ;
        RECT 118.480 199.010 118.765 199.470 ;
        RECT 118.935 198.840 119.205 199.300 ;
        RECT 119.605 199.010 120.005 199.860 ;
        RECT 120.870 199.690 121.320 200.150 ;
        RECT 121.595 199.980 121.875 200.650 ;
        RECT 122.050 200.625 122.505 201.390 ;
        RECT 122.780 201.010 124.080 201.220 ;
        RECT 124.335 201.030 124.665 201.390 ;
        RECT 123.910 200.860 124.080 201.010 ;
        RECT 124.835 200.890 125.095 201.220 ;
        RECT 124.865 200.880 125.095 200.890 ;
        RECT 122.980 200.400 123.200 200.800 ;
        RECT 122.045 200.200 122.535 200.400 ;
        RECT 122.725 200.190 123.200 200.400 ;
        RECT 123.445 200.400 123.655 200.800 ;
        RECT 123.910 200.735 124.665 200.860 ;
        RECT 123.910 200.690 124.755 200.735 ;
        RECT 124.485 200.570 124.755 200.690 ;
        RECT 123.445 200.190 123.775 200.400 ;
        RECT 123.945 200.130 124.355 200.435 ;
        RECT 120.195 199.470 121.320 199.690 ;
        RECT 120.195 199.010 120.475 199.470 ;
        RECT 120.995 198.840 121.320 199.300 ;
        RECT 121.490 199.010 121.875 199.980 ;
        RECT 122.050 199.960 123.225 200.020 ;
        RECT 124.585 199.995 124.755 200.570 ;
        RECT 124.555 199.960 124.755 199.995 ;
        RECT 122.050 199.850 124.755 199.960 ;
        RECT 122.050 199.230 122.305 199.850 ;
        RECT 122.895 199.790 124.695 199.850 ;
        RECT 122.895 199.760 123.225 199.790 ;
        RECT 124.925 199.690 125.095 200.880 ;
        RECT 122.555 199.590 122.740 199.680 ;
        RECT 123.330 199.590 124.165 199.600 ;
        RECT 122.555 199.390 124.165 199.590 ;
        RECT 122.555 199.350 122.785 199.390 ;
        RECT 122.050 199.010 122.385 199.230 ;
        RECT 123.390 198.840 123.745 199.220 ;
        RECT 123.915 199.010 124.165 199.390 ;
        RECT 124.415 198.840 124.665 199.620 ;
        RECT 124.835 199.010 125.095 199.690 ;
        RECT 126.185 200.665 126.445 201.220 ;
        RECT 126.615 200.945 127.045 201.390 ;
        RECT 127.280 200.820 127.450 201.220 ;
        RECT 127.620 200.990 128.340 201.390 ;
        RECT 126.185 199.950 126.360 200.665 ;
        RECT 127.280 200.650 128.160 200.820 ;
        RECT 128.510 200.775 128.680 201.220 ;
        RECT 129.255 200.880 129.655 201.390 ;
        RECT 126.530 200.150 126.785 200.480 ;
        RECT 126.185 199.010 126.445 199.950 ;
        RECT 126.615 199.670 126.785 200.150 ;
        RECT 127.010 199.860 127.340 200.480 ;
        RECT 127.510 200.100 127.800 200.480 ;
        RECT 127.990 199.930 128.160 200.650 ;
        RECT 127.640 199.760 128.160 199.930 ;
        RECT 128.330 200.605 128.680 200.775 ;
        RECT 126.615 199.500 127.375 199.670 ;
        RECT 127.640 199.570 127.810 199.760 ;
        RECT 128.330 199.580 128.500 200.605 ;
        RECT 128.920 200.120 129.180 200.710 ;
        RECT 128.700 199.820 129.180 200.120 ;
        RECT 129.380 199.820 129.640 200.710 ;
        RECT 130.785 200.650 131.170 201.220 ;
        RECT 131.340 200.930 131.665 201.390 ;
        RECT 132.185 200.760 132.465 201.220 ;
        RECT 130.785 199.980 131.065 200.650 ;
        RECT 131.340 200.590 132.465 200.760 ;
        RECT 131.340 200.480 131.790 200.590 ;
        RECT 131.235 200.150 131.790 200.480 ;
        RECT 132.655 200.420 133.055 201.220 ;
        RECT 133.455 200.930 133.725 201.390 ;
        RECT 133.895 200.760 134.180 201.220 ;
        RECT 134.470 200.885 134.805 201.390 ;
        RECT 134.975 200.820 135.215 201.195 ;
        RECT 135.495 201.060 135.665 201.205 ;
        RECT 135.495 200.865 135.870 201.060 ;
        RECT 136.230 200.895 136.625 201.390 ;
        RECT 127.205 199.275 127.375 199.500 ;
        RECT 128.090 199.410 128.500 199.580 ;
        RECT 128.675 199.470 129.615 199.640 ;
        RECT 128.090 199.275 128.345 199.410 ;
        RECT 126.615 198.840 126.945 199.240 ;
        RECT 127.205 199.105 128.345 199.275 ;
        RECT 128.675 199.220 128.845 199.470 ;
        RECT 128.090 199.010 128.345 199.105 ;
        RECT 128.515 199.050 128.845 199.220 ;
        RECT 129.015 198.840 129.265 199.300 ;
        RECT 129.435 199.010 129.615 199.470 ;
        RECT 130.785 199.010 131.170 199.980 ;
        RECT 131.340 199.690 131.790 200.150 ;
        RECT 131.960 199.860 133.055 200.420 ;
        RECT 131.340 199.470 132.465 199.690 ;
        RECT 131.340 198.840 131.665 199.300 ;
        RECT 132.185 199.010 132.465 199.470 ;
        RECT 132.655 199.010 133.055 199.860 ;
        RECT 133.225 200.590 134.180 200.760 ;
        RECT 133.225 199.690 133.435 200.590 ;
        RECT 133.605 199.860 134.295 200.420 ;
        RECT 134.525 199.860 134.825 200.710 ;
        RECT 134.995 200.670 135.215 200.820 ;
        RECT 134.995 200.340 135.530 200.670 ;
        RECT 135.700 200.530 135.870 200.865 ;
        RECT 136.795 200.700 137.035 201.220 ;
        RECT 134.995 199.690 135.230 200.340 ;
        RECT 135.700 200.170 136.685 200.530 ;
        RECT 133.225 199.470 134.180 199.690 ;
        RECT 133.455 198.840 133.725 199.300 ;
        RECT 133.895 199.010 134.180 199.470 ;
        RECT 134.555 199.460 135.230 199.690 ;
        RECT 135.400 200.150 136.685 200.170 ;
        RECT 135.400 200.000 136.260 200.150 ;
        RECT 134.555 199.030 134.725 199.460 ;
        RECT 134.895 198.840 135.225 199.290 ;
        RECT 135.400 199.055 135.685 200.000 ;
        RECT 136.860 199.895 137.035 200.700 ;
        RECT 137.265 200.570 137.495 201.390 ;
        RECT 137.665 200.590 137.995 201.220 ;
        RECT 137.245 200.150 137.575 200.400 ;
        RECT 137.745 199.990 137.995 200.590 ;
        RECT 138.165 200.570 138.375 201.390 ;
        RECT 138.625 200.580 138.865 201.390 ;
        RECT 139.035 200.580 139.365 201.220 ;
        RECT 139.535 200.580 139.805 201.390 ;
        RECT 140.995 200.840 141.165 201.220 ;
        RECT 141.380 201.010 141.710 201.390 ;
        RECT 140.995 200.670 141.710 200.840 ;
        RECT 138.605 200.150 138.955 200.400 ;
        RECT 135.860 199.520 136.555 199.830 ;
        RECT 135.865 198.840 136.550 199.310 ;
        RECT 136.730 199.110 137.035 199.895 ;
        RECT 137.265 198.840 137.495 199.980 ;
        RECT 137.665 199.010 137.995 199.990 ;
        RECT 139.125 199.980 139.295 200.580 ;
        RECT 139.465 200.150 139.815 200.400 ;
        RECT 140.905 200.120 141.260 200.490 ;
        RECT 141.540 200.480 141.710 200.670 ;
        RECT 141.880 200.645 142.135 201.220 ;
        RECT 141.540 200.150 141.795 200.480 ;
        RECT 138.165 198.840 138.375 199.980 ;
        RECT 138.615 199.810 139.295 199.980 ;
        RECT 138.615 199.025 138.945 199.810 ;
        RECT 139.475 198.840 139.805 199.980 ;
        RECT 141.540 199.940 141.710 200.150 ;
        RECT 140.995 199.770 141.710 199.940 ;
        RECT 141.965 199.915 142.135 200.645 ;
        RECT 142.310 200.550 142.570 201.390 ;
        RECT 142.745 200.665 143.035 201.390 ;
        RECT 143.245 200.570 143.475 201.390 ;
        RECT 143.645 200.590 143.975 201.220 ;
        RECT 143.225 200.150 143.555 200.400 ;
        RECT 140.995 199.010 141.165 199.770 ;
        RECT 141.380 198.840 141.710 199.600 ;
        RECT 141.880 199.010 142.135 199.915 ;
        RECT 142.310 198.840 142.570 199.990 ;
        RECT 142.745 198.840 143.035 200.005 ;
        RECT 143.725 199.990 143.975 200.590 ;
        RECT 144.145 200.570 144.355 201.390 ;
        RECT 144.675 200.840 144.845 201.220 ;
        RECT 145.060 201.010 145.390 201.390 ;
        RECT 144.675 200.670 145.390 200.840 ;
        RECT 144.585 200.120 144.940 200.490 ;
        RECT 145.220 200.480 145.390 200.670 ;
        RECT 145.560 200.645 145.815 201.220 ;
        RECT 145.220 200.150 145.475 200.480 ;
        RECT 143.245 198.840 143.475 199.980 ;
        RECT 143.645 199.010 143.975 199.990 ;
        RECT 144.145 198.840 144.355 199.980 ;
        RECT 145.220 199.940 145.390 200.150 ;
        RECT 144.675 199.770 145.390 199.940 ;
        RECT 145.645 199.915 145.815 200.645 ;
        RECT 145.990 200.550 146.250 201.390 ;
        RECT 146.425 200.640 147.635 201.390 ;
        RECT 144.675 199.010 144.845 199.770 ;
        RECT 145.060 198.840 145.390 199.600 ;
        RECT 145.560 199.010 145.815 199.915 ;
        RECT 145.990 198.840 146.250 199.990 ;
        RECT 146.425 199.930 146.945 200.470 ;
        RECT 147.115 200.100 147.635 200.640 ;
        RECT 146.425 198.840 147.635 199.930 ;
        RECT 13.860 198.670 147.720 198.840 ;
        RECT 13.945 197.580 15.155 198.670 ;
        RECT 13.945 196.870 14.465 197.410 ;
        RECT 14.635 197.040 15.155 197.580 ;
        RECT 15.330 197.520 15.590 198.670 ;
        RECT 15.765 197.595 16.020 198.500 ;
        RECT 16.190 197.910 16.520 198.670 ;
        RECT 16.735 197.740 16.905 198.500 ;
        RECT 17.630 198.000 17.885 198.500 ;
        RECT 18.055 198.170 18.385 198.670 ;
        RECT 17.630 197.830 18.380 198.000 ;
        RECT 13.945 196.120 15.155 196.870 ;
        RECT 15.330 196.120 15.590 196.960 ;
        RECT 15.765 196.865 15.935 197.595 ;
        RECT 16.190 197.570 16.905 197.740 ;
        RECT 16.190 197.360 16.360 197.570 ;
        RECT 16.105 197.030 16.360 197.360 ;
        RECT 15.765 196.290 16.020 196.865 ;
        RECT 16.190 196.840 16.360 197.030 ;
        RECT 16.640 197.020 16.995 197.390 ;
        RECT 17.630 197.010 17.980 197.660 ;
        RECT 18.150 196.840 18.380 197.830 ;
        RECT 16.190 196.670 16.905 196.840 ;
        RECT 16.190 196.120 16.520 196.500 ;
        RECT 16.735 196.290 16.905 196.670 ;
        RECT 17.630 196.670 18.380 196.840 ;
        RECT 17.630 196.380 17.885 196.670 ;
        RECT 18.055 196.120 18.385 196.500 ;
        RECT 18.555 196.380 18.725 198.500 ;
        RECT 18.895 197.700 19.220 198.485 ;
        RECT 19.390 198.210 19.640 198.670 ;
        RECT 19.810 198.170 20.060 198.500 ;
        RECT 20.275 198.170 20.955 198.500 ;
        RECT 19.810 198.040 19.980 198.170 ;
        RECT 19.585 197.870 19.980 198.040 ;
        RECT 18.955 196.650 19.415 197.700 ;
        RECT 19.585 196.510 19.755 197.870 ;
        RECT 20.150 197.610 20.615 198.000 ;
        RECT 19.925 196.800 20.275 197.420 ;
        RECT 20.445 197.020 20.615 197.610 ;
        RECT 20.785 197.390 20.955 198.170 ;
        RECT 21.125 198.070 21.295 198.410 ;
        RECT 21.530 198.240 21.860 198.670 ;
        RECT 22.030 198.070 22.200 198.410 ;
        RECT 22.495 198.210 22.865 198.670 ;
        RECT 21.125 197.900 22.200 198.070 ;
        RECT 23.035 198.040 23.205 198.500 ;
        RECT 23.440 198.160 24.310 198.500 ;
        RECT 24.480 198.210 24.730 198.670 ;
        RECT 22.645 197.870 23.205 198.040 ;
        RECT 22.645 197.730 22.815 197.870 ;
        RECT 21.315 197.560 22.815 197.730 ;
        RECT 23.510 197.700 23.970 197.990 ;
        RECT 20.785 197.220 22.475 197.390 ;
        RECT 20.445 196.800 20.800 197.020 ;
        RECT 20.970 196.510 21.140 197.220 ;
        RECT 21.345 196.800 22.135 197.050 ;
        RECT 22.305 197.040 22.475 197.220 ;
        RECT 22.645 196.870 22.815 197.560 ;
        RECT 19.085 196.120 19.415 196.480 ;
        RECT 19.585 196.340 20.080 196.510 ;
        RECT 20.285 196.340 21.140 196.510 ;
        RECT 22.015 196.120 22.345 196.580 ;
        RECT 22.555 196.480 22.815 196.870 ;
        RECT 23.005 197.690 23.970 197.700 ;
        RECT 24.140 197.780 24.310 198.160 ;
        RECT 24.900 198.120 25.070 198.410 ;
        RECT 25.250 198.290 25.580 198.670 ;
        RECT 24.900 197.950 25.700 198.120 ;
        RECT 23.005 197.530 23.680 197.690 ;
        RECT 24.140 197.610 25.360 197.780 ;
        RECT 23.005 196.740 23.215 197.530 ;
        RECT 24.140 197.520 24.310 197.610 ;
        RECT 23.385 196.740 23.735 197.360 ;
        RECT 23.905 197.350 24.310 197.520 ;
        RECT 23.905 196.570 24.075 197.350 ;
        RECT 24.245 196.900 24.465 197.180 ;
        RECT 24.645 197.070 25.185 197.440 ;
        RECT 25.530 197.360 25.700 197.950 ;
        RECT 25.920 197.530 26.225 198.670 ;
        RECT 26.395 197.480 26.650 198.360 ;
        RECT 26.825 197.505 27.115 198.670 ;
        RECT 25.530 197.330 26.270 197.360 ;
        RECT 24.245 196.730 24.775 196.900 ;
        RECT 22.555 196.310 22.905 196.480 ;
        RECT 23.125 196.290 24.075 196.570 ;
        RECT 24.245 196.120 24.435 196.560 ;
        RECT 24.605 196.500 24.775 196.730 ;
        RECT 24.945 196.670 25.185 197.070 ;
        RECT 25.355 197.030 26.270 197.330 ;
        RECT 25.355 196.855 25.680 197.030 ;
        RECT 25.355 196.500 25.675 196.855 ;
        RECT 26.440 196.830 26.650 197.480 ;
        RECT 24.605 196.330 25.675 196.500 ;
        RECT 25.920 196.120 26.225 196.580 ;
        RECT 26.395 196.300 26.650 196.830 ;
        RECT 26.825 196.120 27.115 196.845 ;
        RECT 27.295 196.300 27.555 198.490 ;
        RECT 27.725 197.940 28.065 198.670 ;
        RECT 28.245 197.760 28.515 198.490 ;
        RECT 27.745 197.540 28.515 197.760 ;
        RECT 28.695 197.780 28.925 198.490 ;
        RECT 29.095 197.960 29.425 198.670 ;
        RECT 29.595 197.780 29.855 198.490 ;
        RECT 28.695 197.540 29.855 197.780 ;
        RECT 27.745 196.870 28.035 197.540 ;
        RECT 30.050 197.520 30.310 198.670 ;
        RECT 30.485 197.595 30.740 198.500 ;
        RECT 30.910 197.910 31.240 198.670 ;
        RECT 31.455 197.740 31.625 198.500 ;
        RECT 28.215 197.050 28.680 197.360 ;
        RECT 28.860 197.050 29.385 197.360 ;
        RECT 27.745 196.670 28.975 196.870 ;
        RECT 27.815 196.120 28.485 196.490 ;
        RECT 28.665 196.300 28.975 196.670 ;
        RECT 29.155 196.410 29.385 197.050 ;
        RECT 29.565 197.030 29.865 197.360 ;
        RECT 29.565 196.120 29.855 196.850 ;
        RECT 30.050 196.120 30.310 196.960 ;
        RECT 30.485 196.865 30.655 197.595 ;
        RECT 30.910 197.570 31.625 197.740 ;
        RECT 32.090 197.700 32.420 198.500 ;
        RECT 32.590 197.870 32.920 198.670 ;
        RECT 33.220 197.700 33.550 198.500 ;
        RECT 34.195 197.870 34.445 198.670 ;
        RECT 30.910 197.360 31.080 197.570 ;
        RECT 32.090 197.530 34.525 197.700 ;
        RECT 34.715 197.530 34.885 198.670 ;
        RECT 35.055 197.530 35.395 198.500 ;
        RECT 30.825 197.030 31.080 197.360 ;
        RECT 30.485 196.290 30.740 196.865 ;
        RECT 30.910 196.840 31.080 197.030 ;
        RECT 31.360 197.020 31.715 197.390 ;
        RECT 31.885 197.110 32.235 197.360 ;
        RECT 32.420 196.900 32.590 197.530 ;
        RECT 32.760 197.110 33.090 197.310 ;
        RECT 33.260 197.110 33.590 197.310 ;
        RECT 33.760 197.110 34.180 197.310 ;
        RECT 34.355 197.280 34.525 197.530 ;
        RECT 35.165 197.480 35.395 197.530 ;
        RECT 34.355 197.110 35.050 197.280 ;
        RECT 30.910 196.670 31.625 196.840 ;
        RECT 30.910 196.120 31.240 196.500 ;
        RECT 31.455 196.290 31.625 196.670 ;
        RECT 32.090 196.290 32.590 196.900 ;
        RECT 33.220 196.770 34.445 196.940 ;
        RECT 35.220 196.920 35.395 197.480 ;
        RECT 33.220 196.290 33.550 196.770 ;
        RECT 33.720 196.120 33.945 196.580 ;
        RECT 34.115 196.290 34.445 196.770 ;
        RECT 34.635 196.120 34.885 196.920 ;
        RECT 35.055 196.290 35.395 196.920 ;
        RECT 35.575 196.300 35.835 198.490 ;
        RECT 36.005 197.940 36.345 198.670 ;
        RECT 36.525 197.760 36.795 198.490 ;
        RECT 36.025 197.540 36.795 197.760 ;
        RECT 36.975 197.780 37.205 198.490 ;
        RECT 37.375 197.960 37.705 198.670 ;
        RECT 37.875 197.780 38.135 198.490 ;
        RECT 36.975 197.540 38.135 197.780 ;
        RECT 36.025 196.870 36.315 197.540 ;
        RECT 38.330 197.530 38.605 198.500 ;
        RECT 38.815 197.870 39.095 198.670 ;
        RECT 39.265 198.160 40.455 198.450 ;
        RECT 39.265 197.820 40.435 197.990 ;
        RECT 39.265 197.700 39.435 197.820 ;
        RECT 38.775 197.530 39.435 197.700 ;
        RECT 36.495 197.050 36.960 197.360 ;
        RECT 37.140 197.050 37.665 197.360 ;
        RECT 36.025 196.670 37.255 196.870 ;
        RECT 36.095 196.120 36.765 196.490 ;
        RECT 36.945 196.300 37.255 196.670 ;
        RECT 37.435 196.410 37.665 197.050 ;
        RECT 37.845 197.030 38.145 197.360 ;
        RECT 37.845 196.120 38.135 196.850 ;
        RECT 38.330 196.795 38.500 197.530 ;
        RECT 38.775 197.360 38.945 197.530 ;
        RECT 39.745 197.360 39.940 197.650 ;
        RECT 40.110 197.530 40.435 197.820 ;
        RECT 41.545 197.530 41.825 198.670 ;
        RECT 41.995 197.520 42.325 198.500 ;
        RECT 42.495 197.530 42.755 198.670 ;
        RECT 43.865 197.820 44.195 198.670 ;
        RECT 44.365 198.330 45.475 198.500 ;
        RECT 44.365 197.820 44.585 198.330 ;
        RECT 45.285 198.170 45.475 198.330 ;
        RECT 45.670 198.210 46.000 198.670 ;
        RECT 44.755 198.000 45.055 198.160 ;
        RECT 46.170 198.000 46.405 198.500 ;
        RECT 44.755 197.820 46.405 198.000 ;
        RECT 38.670 197.030 38.945 197.360 ;
        RECT 39.115 197.030 39.940 197.360 ;
        RECT 40.110 197.030 40.455 197.360 ;
        RECT 41.555 197.090 41.890 197.360 ;
        RECT 38.775 196.860 38.945 197.030 ;
        RECT 42.060 196.920 42.230 197.520 ;
        RECT 43.880 197.480 45.855 197.650 ;
        RECT 42.400 197.110 42.735 197.360 ;
        RECT 43.880 197.090 44.210 197.480 ;
        RECT 44.380 197.110 45.180 197.310 ;
        RECT 45.360 197.110 45.855 197.480 ;
        RECT 38.330 196.450 38.605 196.795 ;
        RECT 38.775 196.690 40.440 196.860 ;
        RECT 38.795 196.120 39.175 196.520 ;
        RECT 39.345 196.340 39.515 196.690 ;
        RECT 39.685 196.120 40.015 196.520 ;
        RECT 40.185 196.340 40.440 196.690 ;
        RECT 41.545 196.120 41.855 196.920 ;
        RECT 42.060 196.290 42.755 196.920 ;
        RECT 43.865 196.750 46.025 196.920 ;
        RECT 43.865 196.290 44.195 196.750 ;
        RECT 44.375 196.120 44.545 196.580 ;
        RECT 44.725 196.290 45.055 196.750 ;
        RECT 45.285 196.120 45.455 196.580 ;
        RECT 45.695 196.460 46.025 196.750 ;
        RECT 46.195 196.630 46.405 197.820 ;
        RECT 46.575 197.605 46.885 198.670 ;
        RECT 47.085 197.820 47.415 198.670 ;
        RECT 47.585 198.330 48.695 198.500 ;
        RECT 47.585 197.820 47.805 198.330 ;
        RECT 48.505 198.170 48.695 198.330 ;
        RECT 48.890 198.210 49.220 198.670 ;
        RECT 47.975 198.000 48.275 198.160 ;
        RECT 49.390 198.000 49.625 198.500 ;
        RECT 47.975 197.820 49.625 198.000 ;
        RECT 47.100 197.480 49.135 197.650 ;
        RECT 46.575 196.800 46.890 197.435 ;
        RECT 47.100 197.090 47.430 197.480 ;
        RECT 47.600 197.110 48.400 197.310 ;
        RECT 48.580 197.110 49.075 197.480 ;
        RECT 47.085 196.750 49.245 196.920 ;
        RECT 46.575 196.460 46.885 196.630 ;
        RECT 45.695 196.290 46.885 196.460 ;
        RECT 47.085 196.290 47.415 196.750 ;
        RECT 47.595 196.120 47.765 196.580 ;
        RECT 47.945 196.290 48.275 196.750 ;
        RECT 48.505 196.120 48.675 196.580 ;
        RECT 48.915 196.460 49.245 196.750 ;
        RECT 49.415 196.630 49.625 197.820 ;
        RECT 49.795 197.605 50.105 198.670 ;
        RECT 50.285 197.530 50.545 198.670 ;
        RECT 50.715 197.520 51.045 198.500 ;
        RECT 51.215 197.530 51.495 198.670 ;
        RECT 49.795 196.800 50.110 197.435 ;
        RECT 50.305 197.110 50.640 197.360 ;
        RECT 50.810 196.920 50.980 197.520 ;
        RECT 52.585 197.505 52.875 198.670 ;
        RECT 53.045 197.595 53.315 198.500 ;
        RECT 53.485 197.910 53.815 198.670 ;
        RECT 53.995 197.740 54.165 198.500 ;
        RECT 51.150 197.090 51.485 197.360 ;
        RECT 49.795 196.460 50.105 196.630 ;
        RECT 48.915 196.290 50.105 196.460 ;
        RECT 50.285 196.290 50.980 196.920 ;
        RECT 51.185 196.120 51.495 196.920 ;
        RECT 52.585 196.120 52.875 196.845 ;
        RECT 53.045 196.795 53.215 197.595 ;
        RECT 53.500 197.570 54.165 197.740 ;
        RECT 54.425 197.580 55.635 198.670 ;
        RECT 53.500 197.425 53.670 197.570 ;
        RECT 53.385 197.095 53.670 197.425 ;
        RECT 53.500 196.840 53.670 197.095 ;
        RECT 53.905 197.020 54.235 197.390 ;
        RECT 54.425 196.870 54.945 197.410 ;
        RECT 55.115 197.040 55.635 197.580 ;
        RECT 55.865 197.530 56.075 198.670 ;
        RECT 56.245 197.520 56.575 198.500 ;
        RECT 56.745 197.530 56.975 198.670 ;
        RECT 57.185 197.530 57.465 198.670 ;
        RECT 57.635 197.520 57.965 198.500 ;
        RECT 58.135 197.530 58.395 198.670 ;
        RECT 58.565 197.530 58.825 198.670 ;
        RECT 58.995 197.520 59.325 198.500 ;
        RECT 59.495 197.530 59.775 198.670 ;
        RECT 59.950 198.000 60.205 198.500 ;
        RECT 60.375 198.170 60.705 198.670 ;
        RECT 59.950 197.830 60.700 198.000 ;
        RECT 53.045 196.290 53.305 196.795 ;
        RECT 53.500 196.670 54.165 196.840 ;
        RECT 53.485 196.120 53.815 196.500 ;
        RECT 53.995 196.290 54.165 196.670 ;
        RECT 54.425 196.120 55.635 196.870 ;
        RECT 55.865 196.120 56.075 196.940 ;
        RECT 56.245 196.920 56.495 197.520 ;
        RECT 56.665 197.110 56.995 197.360 ;
        RECT 57.195 197.090 57.530 197.360 ;
        RECT 56.245 196.290 56.575 196.920 ;
        RECT 56.745 196.120 56.975 196.940 ;
        RECT 57.700 196.920 57.870 197.520 ;
        RECT 58.040 197.110 58.375 197.360 ;
        RECT 58.585 197.110 58.920 197.360 ;
        RECT 59.090 196.920 59.260 197.520 ;
        RECT 59.430 197.090 59.765 197.360 ;
        RECT 59.950 197.010 60.300 197.660 ;
        RECT 57.185 196.120 57.495 196.920 ;
        RECT 57.700 196.290 58.395 196.920 ;
        RECT 58.565 196.290 59.260 196.920 ;
        RECT 59.465 196.120 59.775 196.920 ;
        RECT 60.470 196.840 60.700 197.830 ;
        RECT 59.950 196.670 60.700 196.840 ;
        RECT 59.950 196.380 60.205 196.670 ;
        RECT 60.375 196.120 60.705 196.500 ;
        RECT 60.875 196.380 61.045 198.500 ;
        RECT 61.215 197.700 61.540 198.485 ;
        RECT 61.710 198.210 61.960 198.670 ;
        RECT 62.130 198.170 62.380 198.500 ;
        RECT 62.595 198.170 63.275 198.500 ;
        RECT 62.130 198.040 62.300 198.170 ;
        RECT 61.905 197.870 62.300 198.040 ;
        RECT 61.275 196.650 61.735 197.700 ;
        RECT 61.905 196.510 62.075 197.870 ;
        RECT 62.470 197.610 62.935 198.000 ;
        RECT 62.245 196.800 62.595 197.420 ;
        RECT 62.765 197.020 62.935 197.610 ;
        RECT 63.105 197.390 63.275 198.170 ;
        RECT 63.445 198.070 63.615 198.410 ;
        RECT 63.850 198.240 64.180 198.670 ;
        RECT 64.350 198.070 64.520 198.410 ;
        RECT 64.815 198.210 65.185 198.670 ;
        RECT 63.445 197.900 64.520 198.070 ;
        RECT 65.355 198.040 65.525 198.500 ;
        RECT 65.760 198.160 66.630 198.500 ;
        RECT 66.800 198.210 67.050 198.670 ;
        RECT 64.965 197.870 65.525 198.040 ;
        RECT 64.965 197.730 65.135 197.870 ;
        RECT 63.635 197.560 65.135 197.730 ;
        RECT 65.830 197.700 66.290 197.990 ;
        RECT 63.105 197.220 64.795 197.390 ;
        RECT 62.765 196.800 63.120 197.020 ;
        RECT 63.290 196.510 63.460 197.220 ;
        RECT 63.665 196.800 64.455 197.050 ;
        RECT 64.625 197.040 64.795 197.220 ;
        RECT 64.965 196.870 65.135 197.560 ;
        RECT 61.405 196.120 61.735 196.480 ;
        RECT 61.905 196.340 62.400 196.510 ;
        RECT 62.605 196.340 63.460 196.510 ;
        RECT 64.335 196.120 64.665 196.580 ;
        RECT 64.875 196.480 65.135 196.870 ;
        RECT 65.325 197.690 66.290 197.700 ;
        RECT 66.460 197.780 66.630 198.160 ;
        RECT 67.220 198.120 67.390 198.410 ;
        RECT 67.570 198.290 67.900 198.670 ;
        RECT 67.220 197.950 68.020 198.120 ;
        RECT 65.325 197.530 66.000 197.690 ;
        RECT 66.460 197.610 67.680 197.780 ;
        RECT 65.325 196.740 65.535 197.530 ;
        RECT 66.460 197.520 66.630 197.610 ;
        RECT 65.705 196.740 66.055 197.360 ;
        RECT 66.225 197.350 66.630 197.520 ;
        RECT 66.225 196.570 66.395 197.350 ;
        RECT 66.565 196.900 66.785 197.180 ;
        RECT 66.965 197.070 67.505 197.440 ;
        RECT 67.850 197.330 68.020 197.950 ;
        RECT 68.195 197.610 68.365 198.670 ;
        RECT 68.575 197.660 68.865 198.500 ;
        RECT 69.035 197.830 69.205 198.670 ;
        RECT 69.415 197.660 69.665 198.500 ;
        RECT 69.875 197.830 70.045 198.670 ;
        RECT 70.530 198.290 70.865 198.670 ;
        RECT 68.575 197.490 70.300 197.660 ;
        RECT 66.565 196.730 67.095 196.900 ;
        RECT 64.875 196.310 65.225 196.480 ;
        RECT 65.445 196.290 66.395 196.570 ;
        RECT 66.565 196.120 66.755 196.560 ;
        RECT 66.925 196.500 67.095 196.730 ;
        RECT 67.265 196.670 67.505 197.070 ;
        RECT 67.675 197.320 68.020 197.330 ;
        RECT 67.675 197.110 69.705 197.320 ;
        RECT 67.675 196.855 68.000 197.110 ;
        RECT 69.890 196.940 70.300 197.490 ;
        RECT 67.675 196.500 67.995 196.855 ;
        RECT 66.925 196.330 67.995 196.500 ;
        RECT 68.195 196.120 68.365 196.930 ;
        RECT 68.535 196.770 70.300 196.940 ;
        RECT 70.525 196.800 70.765 198.110 ;
        RECT 71.035 197.700 71.285 198.500 ;
        RECT 71.505 197.950 71.835 198.670 ;
        RECT 72.020 197.700 72.270 198.500 ;
        RECT 72.735 197.870 73.065 198.670 ;
        RECT 73.235 198.240 73.575 198.500 ;
        RECT 70.935 197.530 73.125 197.700 ;
        RECT 68.535 196.290 68.865 196.770 ;
        RECT 69.035 196.120 69.205 196.590 ;
        RECT 69.375 196.290 69.705 196.770 ;
        RECT 70.935 196.620 71.105 197.530 ;
        RECT 72.810 197.360 73.125 197.530 ;
        RECT 69.875 196.120 70.045 196.590 ;
        RECT 70.610 196.290 71.105 196.620 ;
        RECT 71.325 196.395 71.675 197.360 ;
        RECT 71.855 196.390 72.155 197.360 ;
        RECT 72.335 196.390 72.615 197.360 ;
        RECT 72.810 197.110 73.140 197.360 ;
        RECT 72.795 196.120 73.065 196.920 ;
        RECT 73.315 196.840 73.575 198.240 ;
        RECT 73.745 198.115 74.350 198.670 ;
        RECT 74.525 198.160 75.005 198.500 ;
        RECT 75.175 198.125 75.430 198.670 ;
        RECT 73.745 198.015 74.360 198.115 ;
        RECT 74.175 197.990 74.360 198.015 ;
        RECT 73.745 197.395 74.005 197.845 ;
        RECT 74.175 197.745 74.505 197.990 ;
        RECT 74.675 197.670 75.430 197.920 ;
        RECT 75.600 197.800 75.875 198.500 ;
        RECT 74.660 197.635 75.430 197.670 ;
        RECT 74.645 197.625 75.430 197.635 ;
        RECT 74.640 197.610 75.535 197.625 ;
        RECT 74.620 197.595 75.535 197.610 ;
        RECT 74.600 197.585 75.535 197.595 ;
        RECT 74.575 197.575 75.535 197.585 ;
        RECT 74.505 197.545 75.535 197.575 ;
        RECT 74.485 197.515 75.535 197.545 ;
        RECT 74.465 197.485 75.535 197.515 ;
        RECT 74.435 197.460 75.535 197.485 ;
        RECT 74.400 197.425 75.535 197.460 ;
        RECT 74.370 197.420 75.535 197.425 ;
        RECT 74.370 197.415 74.760 197.420 ;
        RECT 74.370 197.405 74.735 197.415 ;
        RECT 74.370 197.400 74.720 197.405 ;
        RECT 74.370 197.395 74.705 197.400 ;
        RECT 73.745 197.390 74.705 197.395 ;
        RECT 73.745 197.380 74.695 197.390 ;
        RECT 73.745 197.375 74.685 197.380 ;
        RECT 73.745 197.365 74.675 197.375 ;
        RECT 73.745 197.355 74.670 197.365 ;
        RECT 73.745 197.350 74.665 197.355 ;
        RECT 73.745 197.335 74.655 197.350 ;
        RECT 73.745 197.320 74.650 197.335 ;
        RECT 73.745 197.295 74.640 197.320 ;
        RECT 73.745 197.225 74.635 197.295 ;
        RECT 73.235 196.330 73.575 196.840 ;
        RECT 73.745 196.670 74.295 197.055 ;
        RECT 74.465 196.500 74.635 197.225 ;
        RECT 73.745 196.330 74.635 196.500 ;
        RECT 74.805 196.825 75.135 197.250 ;
        RECT 75.305 197.025 75.535 197.420 ;
        RECT 74.805 196.340 75.025 196.825 ;
        RECT 75.705 196.770 75.875 197.800 ;
        RECT 76.510 197.520 76.770 198.670 ;
        RECT 76.945 197.595 77.200 198.500 ;
        RECT 77.370 197.910 77.700 198.670 ;
        RECT 77.915 197.740 78.085 198.500 ;
        RECT 75.195 196.120 75.445 196.660 ;
        RECT 75.615 196.290 75.875 196.770 ;
        RECT 76.510 196.120 76.770 196.960 ;
        RECT 76.945 196.865 77.115 197.595 ;
        RECT 77.370 197.570 78.085 197.740 ;
        RECT 77.370 197.360 77.540 197.570 ;
        RECT 78.345 197.505 78.635 198.670 ;
        RECT 78.810 198.280 79.145 198.500 ;
        RECT 80.150 198.290 80.505 198.670 ;
        RECT 78.810 197.660 79.065 198.280 ;
        RECT 79.315 198.120 79.545 198.160 ;
        RECT 80.675 198.120 80.925 198.500 ;
        RECT 79.315 197.920 80.925 198.120 ;
        RECT 79.315 197.830 79.500 197.920 ;
        RECT 80.090 197.910 80.925 197.920 ;
        RECT 81.175 197.890 81.425 198.670 ;
        RECT 81.595 197.820 81.855 198.500 ;
        RECT 79.655 197.720 79.985 197.750 ;
        RECT 79.655 197.660 81.455 197.720 ;
        RECT 78.810 197.550 81.515 197.660 ;
        RECT 78.810 197.490 79.985 197.550 ;
        RECT 81.315 197.515 81.515 197.550 ;
        RECT 77.285 197.030 77.540 197.360 ;
        RECT 76.945 196.290 77.200 196.865 ;
        RECT 77.370 196.840 77.540 197.030 ;
        RECT 77.820 197.020 78.175 197.390 ;
        RECT 78.805 197.110 79.295 197.310 ;
        RECT 79.485 197.110 79.960 197.320 ;
        RECT 77.370 196.670 78.085 196.840 ;
        RECT 77.370 196.120 77.700 196.500 ;
        RECT 77.915 196.290 78.085 196.670 ;
        RECT 78.345 196.120 78.635 196.845 ;
        RECT 78.810 196.120 79.265 196.885 ;
        RECT 79.740 196.710 79.960 197.110 ;
        RECT 80.205 197.110 80.535 197.320 ;
        RECT 80.205 196.710 80.415 197.110 ;
        RECT 80.705 197.075 81.115 197.380 ;
        RECT 81.345 196.940 81.515 197.515 ;
        RECT 81.245 196.820 81.515 196.940 ;
        RECT 80.670 196.775 81.515 196.820 ;
        RECT 80.670 196.650 81.425 196.775 ;
        RECT 80.670 196.500 80.840 196.650 ;
        RECT 81.685 196.630 81.855 197.820 ;
        RECT 81.625 196.620 81.855 196.630 ;
        RECT 79.540 196.290 80.840 196.500 ;
        RECT 81.095 196.120 81.425 196.480 ;
        RECT 81.595 196.290 81.855 196.620 ;
        RECT 82.945 197.480 83.405 198.490 ;
        RECT 84.475 198.160 84.805 198.670 ;
        RECT 83.575 197.820 85.535 197.990 ;
        RECT 82.945 196.860 83.115 197.480 ;
        RECT 83.575 197.280 83.745 197.820 ;
        RECT 83.285 197.110 83.745 197.280 ;
        RECT 83.925 197.030 84.165 197.650 ;
        RECT 84.335 197.030 84.675 197.650 ;
        RECT 84.845 197.030 85.195 197.650 ;
        RECT 85.365 196.860 85.535 197.820 ;
        RECT 85.705 197.580 89.215 198.670 ;
        RECT 89.385 197.580 90.595 198.670 ;
        RECT 82.945 196.690 84.305 196.860 ;
        RECT 82.945 196.290 83.465 196.690 ;
        RECT 83.635 196.120 83.965 196.520 ;
        RECT 84.135 196.345 84.305 196.690 ;
        RECT 84.475 196.120 84.805 196.860 ;
        RECT 85.040 196.690 85.535 196.860 ;
        RECT 85.705 196.890 87.355 197.410 ;
        RECT 87.525 197.060 89.215 197.580 ;
        RECT 85.040 196.440 85.210 196.690 ;
        RECT 85.705 196.120 89.215 196.890 ;
        RECT 89.385 196.870 89.905 197.410 ;
        RECT 90.075 197.040 90.595 197.580 ;
        RECT 90.775 197.530 91.105 198.670 ;
        RECT 91.635 197.700 91.965 198.485 ;
        RECT 92.145 198.235 97.490 198.670 ;
        RECT 98.130 198.290 98.465 198.670 ;
        RECT 91.285 197.530 91.965 197.700 ;
        RECT 90.765 197.110 91.115 197.360 ;
        RECT 91.285 196.930 91.455 197.530 ;
        RECT 91.625 197.110 91.975 197.360 ;
        RECT 89.385 196.120 90.595 196.870 ;
        RECT 90.775 196.120 91.045 196.930 ;
        RECT 91.215 196.290 91.545 196.930 ;
        RECT 91.715 196.120 91.955 196.930 ;
        RECT 93.730 196.665 94.070 197.495 ;
        RECT 95.550 196.985 95.900 198.235 ;
        RECT 98.125 196.800 98.365 198.110 ;
        RECT 98.635 197.700 98.885 198.500 ;
        RECT 99.105 197.950 99.435 198.670 ;
        RECT 99.620 197.700 99.870 198.500 ;
        RECT 100.335 197.870 100.665 198.670 ;
        RECT 100.835 198.240 101.175 198.500 ;
        RECT 98.535 197.530 100.725 197.700 ;
        RECT 92.145 196.120 97.490 196.665 ;
        RECT 98.535 196.620 98.705 197.530 ;
        RECT 100.410 197.360 100.725 197.530 ;
        RECT 98.210 196.290 98.705 196.620 ;
        RECT 98.925 196.395 99.275 197.360 ;
        RECT 99.455 196.390 99.755 197.360 ;
        RECT 99.935 196.390 100.215 197.360 ;
        RECT 100.410 197.110 100.740 197.360 ;
        RECT 100.395 196.120 100.665 196.920 ;
        RECT 100.915 196.840 101.175 198.240 ;
        RECT 102.075 198.160 102.405 198.670 ;
        RECT 100.835 196.330 101.175 196.840 ;
        RECT 101.345 197.820 103.305 197.990 ;
        RECT 101.345 196.860 101.515 197.820 ;
        RECT 101.685 197.030 102.035 197.650 ;
        RECT 102.205 197.030 102.545 197.650 ;
        RECT 102.715 197.030 102.955 197.650 ;
        RECT 103.135 197.280 103.305 197.820 ;
        RECT 103.475 197.480 103.935 198.490 ;
        RECT 104.105 197.505 104.395 198.670 ;
        RECT 104.570 198.290 104.905 198.670 ;
        RECT 103.135 197.110 103.595 197.280 ;
        RECT 103.765 196.860 103.935 197.480 ;
        RECT 101.345 196.690 101.840 196.860 ;
        RECT 101.670 196.440 101.840 196.690 ;
        RECT 102.075 196.120 102.405 196.860 ;
        RECT 102.575 196.690 103.935 196.860 ;
        RECT 102.575 196.345 102.745 196.690 ;
        RECT 102.915 196.120 103.245 196.520 ;
        RECT 103.415 196.290 103.935 196.690 ;
        RECT 104.105 196.120 104.395 196.845 ;
        RECT 104.565 196.800 104.805 198.110 ;
        RECT 105.075 197.700 105.325 198.500 ;
        RECT 105.545 197.950 105.875 198.670 ;
        RECT 106.060 197.700 106.310 198.500 ;
        RECT 106.775 197.870 107.105 198.670 ;
        RECT 107.275 198.240 107.615 198.500 ;
        RECT 104.975 197.530 107.165 197.700 ;
        RECT 104.975 196.620 105.145 197.530 ;
        RECT 106.850 197.360 107.165 197.530 ;
        RECT 104.650 196.290 105.145 196.620 ;
        RECT 105.365 196.395 105.715 197.360 ;
        RECT 105.895 196.390 106.195 197.360 ;
        RECT 106.375 196.390 106.655 197.360 ;
        RECT 106.850 197.110 107.180 197.360 ;
        RECT 106.835 196.120 107.105 196.920 ;
        RECT 107.355 196.840 107.615 198.240 ;
        RECT 107.785 198.160 108.045 198.670 ;
        RECT 107.785 197.110 108.125 197.990 ;
        RECT 108.295 197.280 108.465 198.500 ;
        RECT 108.705 198.165 109.320 198.670 ;
        RECT 108.705 197.630 108.955 197.995 ;
        RECT 109.125 197.990 109.320 198.165 ;
        RECT 109.490 198.160 109.965 198.500 ;
        RECT 110.135 198.125 110.350 198.670 ;
        RECT 109.125 197.800 109.455 197.990 ;
        RECT 109.675 197.630 110.390 197.925 ;
        RECT 110.560 197.800 110.835 198.500 ;
        RECT 111.010 198.000 111.265 198.500 ;
        RECT 111.435 198.170 111.765 198.670 ;
        RECT 111.010 197.830 111.760 198.000 ;
        RECT 108.705 197.460 110.495 197.630 ;
        RECT 108.295 197.030 109.090 197.280 ;
        RECT 108.295 196.940 108.545 197.030 ;
        RECT 107.275 196.330 107.615 196.840 ;
        RECT 107.785 196.120 108.045 196.940 ;
        RECT 108.215 196.520 108.545 196.940 ;
        RECT 109.260 196.605 109.515 197.460 ;
        RECT 108.725 196.340 109.515 196.605 ;
        RECT 109.685 196.760 110.095 197.280 ;
        RECT 110.265 197.030 110.495 197.460 ;
        RECT 110.665 196.770 110.835 197.800 ;
        RECT 111.010 197.010 111.360 197.660 ;
        RECT 111.530 196.840 111.760 197.830 ;
        RECT 109.685 196.340 109.885 196.760 ;
        RECT 110.075 196.120 110.405 196.580 ;
        RECT 110.575 196.290 110.835 196.770 ;
        RECT 111.010 196.670 111.760 196.840 ;
        RECT 111.010 196.380 111.265 196.670 ;
        RECT 111.435 196.120 111.765 196.500 ;
        RECT 111.935 196.380 112.105 198.500 ;
        RECT 112.275 197.700 112.600 198.485 ;
        RECT 112.770 198.210 113.020 198.670 ;
        RECT 113.190 198.170 113.440 198.500 ;
        RECT 113.655 198.170 114.335 198.500 ;
        RECT 113.190 198.040 113.360 198.170 ;
        RECT 112.965 197.870 113.360 198.040 ;
        RECT 112.335 196.650 112.795 197.700 ;
        RECT 112.965 196.510 113.135 197.870 ;
        RECT 113.530 197.610 113.995 198.000 ;
        RECT 113.305 196.800 113.655 197.420 ;
        RECT 113.825 197.020 113.995 197.610 ;
        RECT 114.165 197.390 114.335 198.170 ;
        RECT 114.505 198.070 114.675 198.410 ;
        RECT 114.910 198.240 115.240 198.670 ;
        RECT 115.410 198.070 115.580 198.410 ;
        RECT 115.875 198.210 116.245 198.670 ;
        RECT 114.505 197.900 115.580 198.070 ;
        RECT 116.415 198.040 116.585 198.500 ;
        RECT 116.820 198.160 117.690 198.500 ;
        RECT 117.860 198.210 118.110 198.670 ;
        RECT 116.025 197.870 116.585 198.040 ;
        RECT 116.025 197.730 116.195 197.870 ;
        RECT 114.695 197.560 116.195 197.730 ;
        RECT 116.890 197.700 117.350 197.990 ;
        RECT 114.165 197.220 115.855 197.390 ;
        RECT 113.825 196.800 114.180 197.020 ;
        RECT 114.350 196.510 114.520 197.220 ;
        RECT 114.725 196.800 115.515 197.050 ;
        RECT 115.685 197.040 115.855 197.220 ;
        RECT 116.025 196.870 116.195 197.560 ;
        RECT 112.465 196.120 112.795 196.480 ;
        RECT 112.965 196.340 113.460 196.510 ;
        RECT 113.665 196.340 114.520 196.510 ;
        RECT 115.395 196.120 115.725 196.580 ;
        RECT 115.935 196.480 116.195 196.870 ;
        RECT 116.385 197.690 117.350 197.700 ;
        RECT 117.520 197.780 117.690 198.160 ;
        RECT 118.280 198.120 118.450 198.410 ;
        RECT 118.630 198.290 118.960 198.670 ;
        RECT 118.280 197.950 119.080 198.120 ;
        RECT 116.385 197.530 117.060 197.690 ;
        RECT 117.520 197.610 118.740 197.780 ;
        RECT 116.385 196.740 116.595 197.530 ;
        RECT 117.520 197.520 117.690 197.610 ;
        RECT 116.765 196.740 117.115 197.360 ;
        RECT 117.285 197.350 117.690 197.520 ;
        RECT 117.285 196.570 117.455 197.350 ;
        RECT 117.625 196.900 117.845 197.180 ;
        RECT 118.025 197.070 118.565 197.440 ;
        RECT 118.910 197.330 119.080 197.950 ;
        RECT 119.255 197.610 119.425 198.670 ;
        RECT 119.635 197.660 119.925 198.500 ;
        RECT 120.095 197.830 120.265 198.670 ;
        RECT 120.475 197.660 120.725 198.500 ;
        RECT 120.935 197.830 121.105 198.670 ;
        RECT 119.635 197.490 121.360 197.660 ;
        RECT 117.625 196.730 118.155 196.900 ;
        RECT 115.935 196.310 116.285 196.480 ;
        RECT 116.505 196.290 117.455 196.570 ;
        RECT 117.625 196.120 117.815 196.560 ;
        RECT 117.985 196.500 118.155 196.730 ;
        RECT 118.325 196.670 118.565 197.070 ;
        RECT 118.735 197.320 119.080 197.330 ;
        RECT 118.735 197.110 120.765 197.320 ;
        RECT 118.735 196.855 119.060 197.110 ;
        RECT 120.950 196.940 121.360 197.490 ;
        RECT 118.735 196.500 119.055 196.855 ;
        RECT 117.985 196.330 119.055 196.500 ;
        RECT 119.255 196.120 119.425 196.930 ;
        RECT 119.595 196.770 121.360 196.940 ;
        RECT 121.585 197.530 121.970 198.500 ;
        RECT 122.140 198.210 122.465 198.670 ;
        RECT 122.985 198.040 123.265 198.500 ;
        RECT 122.140 197.820 123.265 198.040 ;
        RECT 121.585 196.860 121.865 197.530 ;
        RECT 122.140 197.360 122.590 197.820 ;
        RECT 123.455 197.650 123.855 198.500 ;
        RECT 124.255 198.210 124.525 198.670 ;
        RECT 124.695 198.040 124.980 198.500 ;
        RECT 122.035 197.030 122.590 197.360 ;
        RECT 122.760 197.090 123.855 197.650 ;
        RECT 122.140 196.920 122.590 197.030 ;
        RECT 119.595 196.290 119.925 196.770 ;
        RECT 120.095 196.120 120.265 196.590 ;
        RECT 120.435 196.290 120.765 196.770 ;
        RECT 120.935 196.120 121.105 196.590 ;
        RECT 121.585 196.290 121.970 196.860 ;
        RECT 122.140 196.750 123.265 196.920 ;
        RECT 122.140 196.120 122.465 196.580 ;
        RECT 122.985 196.290 123.265 196.750 ;
        RECT 123.455 196.290 123.855 197.090 ;
        RECT 124.025 197.820 124.980 198.040 ;
        RECT 125.275 197.950 125.605 198.670 ;
        RECT 124.025 196.920 124.235 197.820 ;
        RECT 124.405 197.090 125.095 197.650 ;
        RECT 125.265 197.310 125.495 197.650 ;
        RECT 125.785 197.310 126.000 198.425 ;
        RECT 126.195 197.725 126.525 198.500 ;
        RECT 126.695 197.895 127.405 198.670 ;
        RECT 126.195 197.510 127.345 197.725 ;
        RECT 125.265 197.110 125.595 197.310 ;
        RECT 125.785 197.130 126.235 197.310 ;
        RECT 125.905 197.110 126.235 197.130 ;
        RECT 126.405 197.110 126.875 197.340 ;
        RECT 127.060 196.940 127.345 197.510 ;
        RECT 127.575 197.065 127.855 198.500 ;
        RECT 128.030 197.520 128.290 198.670 ;
        RECT 128.465 197.595 128.720 198.500 ;
        RECT 128.890 197.910 129.220 198.670 ;
        RECT 129.435 197.740 129.605 198.500 ;
        RECT 124.025 196.750 124.980 196.920 ;
        RECT 124.255 196.120 124.525 196.580 ;
        RECT 124.695 196.290 124.980 196.750 ;
        RECT 125.265 196.750 126.445 196.940 ;
        RECT 125.265 196.290 125.605 196.750 ;
        RECT 126.115 196.670 126.445 196.750 ;
        RECT 126.635 196.750 127.345 196.940 ;
        RECT 126.635 196.610 126.935 196.750 ;
        RECT 126.620 196.600 126.935 196.610 ;
        RECT 126.610 196.590 126.935 196.600 ;
        RECT 126.600 196.585 126.935 196.590 ;
        RECT 125.775 196.120 125.945 196.580 ;
        RECT 126.595 196.575 126.935 196.585 ;
        RECT 126.590 196.570 126.935 196.575 ;
        RECT 126.585 196.560 126.935 196.570 ;
        RECT 126.580 196.555 126.935 196.560 ;
        RECT 126.575 196.290 126.935 196.555 ;
        RECT 127.175 196.120 127.345 196.580 ;
        RECT 127.515 196.290 127.855 197.065 ;
        RECT 128.030 196.120 128.290 196.960 ;
        RECT 128.465 196.865 128.635 197.595 ;
        RECT 128.890 197.570 129.605 197.740 ;
        RECT 128.890 197.360 129.060 197.570 ;
        RECT 129.865 197.505 130.155 198.670 ;
        RECT 131.305 198.320 133.375 198.490 ;
        RECT 131.305 197.820 131.565 198.320 ;
        RECT 132.235 198.290 133.375 198.320 ;
        RECT 131.735 197.820 132.065 198.140 ;
        RECT 132.235 197.820 132.425 198.290 ;
        RECT 128.805 197.030 129.060 197.360 ;
        RECT 128.465 196.290 128.720 196.865 ;
        RECT 128.890 196.840 129.060 197.030 ;
        RECT 129.340 197.020 129.695 197.390 ;
        RECT 131.260 197.030 131.565 197.650 ;
        RECT 131.735 196.890 132.015 197.820 ;
        RECT 132.595 197.690 132.925 198.110 ;
        RECT 133.095 197.870 133.375 198.290 ;
        RECT 133.595 197.870 133.825 198.670 ;
        RECT 134.005 197.690 134.275 198.500 ;
        RECT 134.455 197.870 134.685 198.670 ;
        RECT 134.865 197.690 135.135 198.500 ;
        RECT 135.315 197.870 135.545 198.670 ;
        RECT 132.195 197.320 132.415 197.650 ;
        RECT 132.595 197.490 135.135 197.690 ;
        RECT 135.335 197.320 135.660 197.690 ;
        RECT 132.195 197.070 132.945 197.320 ;
        RECT 133.530 197.070 134.240 197.320 ;
        RECT 134.900 197.070 135.660 197.320 ;
        RECT 135.845 197.595 136.115 198.500 ;
        RECT 136.285 197.910 136.615 198.670 ;
        RECT 136.795 197.740 136.965 198.500 ;
        RECT 128.890 196.670 129.605 196.840 ;
        RECT 128.890 196.120 129.220 196.500 ;
        RECT 129.435 196.290 129.605 196.670 ;
        RECT 129.865 196.120 130.155 196.845 ;
        RECT 131.305 196.120 131.555 196.850 ;
        RECT 131.735 196.690 134.305 196.890 ;
        RECT 131.735 196.290 131.995 196.690 ;
        RECT 132.165 196.120 132.495 196.510 ;
        RECT 132.665 196.320 132.855 196.690 ;
        RECT 134.485 196.670 135.595 196.890 ;
        RECT 134.485 196.510 134.655 196.670 ;
        RECT 133.025 196.120 133.355 196.510 ;
        RECT 133.545 196.300 134.655 196.510 ;
        RECT 134.835 196.120 135.165 196.490 ;
        RECT 135.345 196.300 135.595 196.670 ;
        RECT 135.845 196.795 136.015 197.595 ;
        RECT 136.300 197.570 136.965 197.740 ;
        RECT 137.315 197.740 137.485 198.500 ;
        RECT 137.700 197.910 138.030 198.670 ;
        RECT 137.315 197.570 138.030 197.740 ;
        RECT 138.200 197.595 138.455 198.500 ;
        RECT 136.300 197.425 136.470 197.570 ;
        RECT 136.185 197.095 136.470 197.425 ;
        RECT 136.300 196.840 136.470 197.095 ;
        RECT 136.705 197.020 137.035 197.390 ;
        RECT 137.225 197.020 137.580 197.390 ;
        RECT 137.860 197.360 138.030 197.570 ;
        RECT 137.860 197.030 138.115 197.360 ;
        RECT 137.860 196.840 138.030 197.030 ;
        RECT 138.285 196.865 138.455 197.595 ;
        RECT 138.630 197.520 138.890 198.670 ;
        RECT 139.155 197.740 139.325 198.500 ;
        RECT 139.540 197.910 139.870 198.670 ;
        RECT 139.155 197.570 139.870 197.740 ;
        RECT 140.040 197.595 140.295 198.500 ;
        RECT 139.065 197.020 139.420 197.390 ;
        RECT 139.700 197.360 139.870 197.570 ;
        RECT 139.700 197.030 139.955 197.360 ;
        RECT 135.845 196.290 136.105 196.795 ;
        RECT 136.300 196.670 136.965 196.840 ;
        RECT 136.285 196.120 136.615 196.500 ;
        RECT 136.795 196.290 136.965 196.670 ;
        RECT 137.315 196.670 138.030 196.840 ;
        RECT 137.315 196.290 137.485 196.670 ;
        RECT 137.700 196.120 138.030 196.500 ;
        RECT 138.200 196.290 138.455 196.865 ;
        RECT 138.630 196.120 138.890 196.960 ;
        RECT 139.700 196.840 139.870 197.030 ;
        RECT 140.125 196.865 140.295 197.595 ;
        RECT 140.470 197.520 140.730 198.670 ;
        RECT 140.995 197.740 141.165 198.500 ;
        RECT 141.380 197.910 141.710 198.670 ;
        RECT 140.995 197.570 141.710 197.740 ;
        RECT 141.880 197.595 142.135 198.500 ;
        RECT 140.905 197.020 141.260 197.390 ;
        RECT 141.540 197.360 141.710 197.570 ;
        RECT 141.540 197.030 141.795 197.360 ;
        RECT 139.155 196.670 139.870 196.840 ;
        RECT 139.155 196.290 139.325 196.670 ;
        RECT 139.540 196.120 139.870 196.500 ;
        RECT 140.040 196.290 140.295 196.865 ;
        RECT 140.470 196.120 140.730 196.960 ;
        RECT 141.540 196.840 141.710 197.030 ;
        RECT 141.965 196.865 142.135 197.595 ;
        RECT 142.310 197.520 142.570 198.670 ;
        RECT 142.835 197.740 143.005 198.500 ;
        RECT 143.220 197.910 143.550 198.670 ;
        RECT 142.835 197.570 143.550 197.740 ;
        RECT 143.720 197.595 143.975 198.500 ;
        RECT 142.745 197.020 143.100 197.390 ;
        RECT 143.380 197.360 143.550 197.570 ;
        RECT 143.380 197.030 143.635 197.360 ;
        RECT 140.995 196.670 141.710 196.840 ;
        RECT 140.995 196.290 141.165 196.670 ;
        RECT 141.380 196.120 141.710 196.500 ;
        RECT 141.880 196.290 142.135 196.865 ;
        RECT 142.310 196.120 142.570 196.960 ;
        RECT 143.380 196.840 143.550 197.030 ;
        RECT 143.805 196.865 143.975 197.595 ;
        RECT 144.150 197.520 144.410 198.670 ;
        RECT 144.675 197.740 144.845 198.500 ;
        RECT 145.060 197.910 145.390 198.670 ;
        RECT 144.675 197.570 145.390 197.740 ;
        RECT 145.560 197.595 145.815 198.500 ;
        RECT 144.585 197.020 144.940 197.390 ;
        RECT 145.220 197.360 145.390 197.570 ;
        RECT 145.220 197.030 145.475 197.360 ;
        RECT 142.835 196.670 143.550 196.840 ;
        RECT 142.835 196.290 143.005 196.670 ;
        RECT 143.220 196.120 143.550 196.500 ;
        RECT 143.720 196.290 143.975 196.865 ;
        RECT 144.150 196.120 144.410 196.960 ;
        RECT 145.220 196.840 145.390 197.030 ;
        RECT 145.645 196.865 145.815 197.595 ;
        RECT 145.990 197.520 146.250 198.670 ;
        RECT 146.425 197.580 147.635 198.670 ;
        RECT 146.425 197.040 146.945 197.580 ;
        RECT 144.675 196.670 145.390 196.840 ;
        RECT 144.675 196.290 144.845 196.670 ;
        RECT 145.060 196.120 145.390 196.500 ;
        RECT 145.560 196.290 145.815 196.865 ;
        RECT 145.990 196.120 146.250 196.960 ;
        RECT 147.115 196.870 147.635 197.410 ;
        RECT 146.425 196.120 147.635 196.870 ;
        RECT 13.860 195.950 147.720 196.120 ;
        RECT 13.945 195.200 15.155 195.950 ;
        RECT 13.945 194.660 14.465 195.200 ;
        RECT 15.330 195.110 15.590 195.950 ;
        RECT 15.765 195.205 16.020 195.780 ;
        RECT 16.190 195.570 16.520 195.950 ;
        RECT 16.735 195.400 16.905 195.780 ;
        RECT 16.190 195.230 16.905 195.400 ;
        RECT 14.635 194.490 15.155 195.030 ;
        RECT 13.945 193.400 15.155 194.490 ;
        RECT 15.330 193.400 15.590 194.550 ;
        RECT 15.765 194.475 15.935 195.205 ;
        RECT 16.190 195.040 16.360 195.230 ;
        RECT 17.170 195.110 17.430 195.950 ;
        RECT 17.605 195.205 17.860 195.780 ;
        RECT 18.030 195.570 18.360 195.950 ;
        RECT 18.575 195.400 18.745 195.780 ;
        RECT 18.030 195.230 18.745 195.400 ;
        RECT 19.010 195.400 19.265 195.690 ;
        RECT 19.435 195.570 19.765 195.950 ;
        RECT 19.010 195.230 19.760 195.400 ;
        RECT 16.105 194.710 16.360 195.040 ;
        RECT 16.190 194.500 16.360 194.710 ;
        RECT 16.640 194.680 16.995 195.050 ;
        RECT 15.765 193.570 16.020 194.475 ;
        RECT 16.190 194.330 16.905 194.500 ;
        RECT 16.190 193.400 16.520 194.160 ;
        RECT 16.735 193.570 16.905 194.330 ;
        RECT 17.170 193.400 17.430 194.550 ;
        RECT 17.605 194.475 17.775 195.205 ;
        RECT 18.030 195.040 18.200 195.230 ;
        RECT 17.945 194.710 18.200 195.040 ;
        RECT 18.030 194.500 18.200 194.710 ;
        RECT 18.480 194.680 18.835 195.050 ;
        RECT 17.605 193.570 17.860 194.475 ;
        RECT 18.030 194.330 18.745 194.500 ;
        RECT 19.010 194.410 19.360 195.060 ;
        RECT 18.030 193.400 18.360 194.160 ;
        RECT 18.575 193.570 18.745 194.330 ;
        RECT 19.530 194.240 19.760 195.230 ;
        RECT 19.010 194.070 19.760 194.240 ;
        RECT 19.010 193.570 19.265 194.070 ;
        RECT 19.435 193.400 19.765 193.900 ;
        RECT 19.935 193.570 20.105 195.690 ;
        RECT 20.465 195.590 20.795 195.950 ;
        RECT 20.965 195.560 21.460 195.730 ;
        RECT 21.665 195.560 22.520 195.730 ;
        RECT 20.335 194.370 20.795 195.420 ;
        RECT 20.275 193.585 20.600 194.370 ;
        RECT 20.965 194.200 21.135 195.560 ;
        RECT 21.305 194.650 21.655 195.270 ;
        RECT 21.825 195.050 22.180 195.270 ;
        RECT 21.825 194.460 21.995 195.050 ;
        RECT 22.350 194.850 22.520 195.560 ;
        RECT 23.395 195.490 23.725 195.950 ;
        RECT 23.935 195.590 24.285 195.760 ;
        RECT 22.725 195.020 23.515 195.270 ;
        RECT 23.935 195.200 24.195 195.590 ;
        RECT 24.505 195.500 25.455 195.780 ;
        RECT 25.625 195.510 25.815 195.950 ;
        RECT 25.985 195.570 27.055 195.740 ;
        RECT 23.685 194.850 23.855 195.030 ;
        RECT 20.965 194.030 21.360 194.200 ;
        RECT 21.530 194.070 21.995 194.460 ;
        RECT 22.165 194.680 23.855 194.850 ;
        RECT 21.190 193.900 21.360 194.030 ;
        RECT 22.165 193.900 22.335 194.680 ;
        RECT 24.025 194.510 24.195 195.200 ;
        RECT 22.695 194.340 24.195 194.510 ;
        RECT 24.385 194.540 24.595 195.330 ;
        RECT 24.765 194.710 25.115 195.330 ;
        RECT 25.285 194.720 25.455 195.500 ;
        RECT 25.985 195.340 26.155 195.570 ;
        RECT 25.625 195.170 26.155 195.340 ;
        RECT 25.625 194.890 25.845 195.170 ;
        RECT 26.325 195.000 26.565 195.400 ;
        RECT 25.285 194.550 25.690 194.720 ;
        RECT 26.025 194.630 26.565 195.000 ;
        RECT 26.735 195.215 27.055 195.570 ;
        RECT 26.735 194.960 27.060 195.215 ;
        RECT 27.255 195.140 27.425 195.950 ;
        RECT 27.595 195.300 27.925 195.780 ;
        RECT 28.095 195.480 28.265 195.950 ;
        RECT 28.435 195.300 28.765 195.780 ;
        RECT 28.935 195.480 29.105 195.950 ;
        RECT 29.585 195.450 29.845 195.780 ;
        RECT 30.015 195.590 30.345 195.950 ;
        RECT 30.600 195.570 31.900 195.780 ;
        RECT 29.585 195.440 29.815 195.450 ;
        RECT 27.595 195.130 29.360 195.300 ;
        RECT 26.735 194.750 28.765 194.960 ;
        RECT 26.735 194.740 27.080 194.750 ;
        RECT 24.385 194.380 25.060 194.540 ;
        RECT 25.520 194.460 25.690 194.550 ;
        RECT 24.385 194.370 25.350 194.380 ;
        RECT 24.025 194.200 24.195 194.340 ;
        RECT 20.770 193.400 21.020 193.860 ;
        RECT 21.190 193.570 21.440 193.900 ;
        RECT 21.655 193.570 22.335 193.900 ;
        RECT 22.505 194.000 23.580 194.170 ;
        RECT 24.025 194.030 24.585 194.200 ;
        RECT 24.890 194.080 25.350 194.370 ;
        RECT 25.520 194.290 26.740 194.460 ;
        RECT 22.505 193.660 22.675 194.000 ;
        RECT 22.910 193.400 23.240 193.830 ;
        RECT 23.410 193.660 23.580 194.000 ;
        RECT 23.875 193.400 24.245 193.860 ;
        RECT 24.415 193.570 24.585 194.030 ;
        RECT 25.520 193.910 25.690 194.290 ;
        RECT 26.910 194.120 27.080 194.740 ;
        RECT 28.950 194.580 29.360 195.130 ;
        RECT 24.820 193.570 25.690 193.910 ;
        RECT 26.280 193.950 27.080 194.120 ;
        RECT 25.860 193.400 26.110 193.860 ;
        RECT 26.280 193.660 26.450 193.950 ;
        RECT 26.630 193.400 26.960 193.780 ;
        RECT 27.255 193.400 27.425 194.460 ;
        RECT 27.635 194.410 29.360 194.580 ;
        RECT 27.635 193.570 27.925 194.410 ;
        RECT 28.095 193.400 28.265 194.240 ;
        RECT 28.475 193.570 28.725 194.410 ;
        RECT 29.585 194.250 29.755 195.440 ;
        RECT 30.600 195.420 30.770 195.570 ;
        RECT 30.015 195.295 30.770 195.420 ;
        RECT 29.925 195.250 30.770 195.295 ;
        RECT 29.925 195.130 30.195 195.250 ;
        RECT 29.925 194.555 30.095 195.130 ;
        RECT 30.325 194.690 30.735 194.995 ;
        RECT 31.025 194.960 31.235 195.360 ;
        RECT 30.905 194.750 31.235 194.960 ;
        RECT 31.480 194.960 31.700 195.360 ;
        RECT 32.175 195.185 32.630 195.950 ;
        RECT 32.805 195.130 33.065 195.950 ;
        RECT 33.235 195.130 33.565 195.550 ;
        RECT 33.745 195.380 34.005 195.780 ;
        RECT 34.175 195.550 34.505 195.950 ;
        RECT 34.675 195.380 34.845 195.730 ;
        RECT 35.015 195.550 35.390 195.950 ;
        RECT 33.745 195.210 35.410 195.380 ;
        RECT 35.580 195.275 35.855 195.620 ;
        RECT 33.315 195.040 33.565 195.130 ;
        RECT 35.240 195.040 35.410 195.210 ;
        RECT 31.480 194.750 31.955 194.960 ;
        RECT 32.145 194.760 32.635 194.960 ;
        RECT 32.810 194.710 33.145 194.960 ;
        RECT 33.315 194.710 34.030 195.040 ;
        RECT 34.245 194.710 35.070 195.040 ;
        RECT 35.240 194.710 35.515 195.040 ;
        RECT 29.925 194.520 30.125 194.555 ;
        RECT 31.455 194.520 32.630 194.580 ;
        RECT 29.925 194.410 32.630 194.520 ;
        RECT 29.985 194.350 31.785 194.410 ;
        RECT 31.455 194.320 31.785 194.350 ;
        RECT 28.935 193.400 29.105 194.240 ;
        RECT 29.585 193.570 29.845 194.250 ;
        RECT 30.015 193.400 30.265 194.180 ;
        RECT 30.515 194.150 31.350 194.160 ;
        RECT 31.940 194.150 32.125 194.240 ;
        RECT 30.515 193.950 32.125 194.150 ;
        RECT 30.515 193.570 30.765 193.950 ;
        RECT 31.895 193.910 32.125 193.950 ;
        RECT 32.375 193.790 32.630 194.410 ;
        RECT 30.935 193.400 31.290 193.780 ;
        RECT 32.295 193.570 32.630 193.790 ;
        RECT 32.805 193.400 33.065 194.540 ;
        RECT 33.315 194.150 33.485 194.710 ;
        RECT 33.745 194.250 34.075 194.540 ;
        RECT 34.245 194.420 34.490 194.710 ;
        RECT 35.240 194.540 35.410 194.710 ;
        RECT 35.685 194.540 35.855 195.275 ;
        RECT 36.525 195.130 36.755 195.950 ;
        RECT 36.925 195.150 37.255 195.780 ;
        RECT 36.505 194.710 36.835 194.960 ;
        RECT 37.005 194.550 37.255 195.150 ;
        RECT 37.425 195.130 37.635 195.950 ;
        RECT 37.935 195.550 38.265 195.950 ;
        RECT 38.435 195.380 38.605 195.650 ;
        RECT 38.775 195.550 39.105 195.950 ;
        RECT 39.275 195.380 39.530 195.650 ;
        RECT 34.750 194.370 35.410 194.540 ;
        RECT 34.750 194.250 34.920 194.370 ;
        RECT 33.745 194.080 34.920 194.250 ;
        RECT 33.305 193.580 34.920 193.910 ;
        RECT 35.090 193.400 35.370 194.200 ;
        RECT 35.580 193.570 35.855 194.540 ;
        RECT 36.525 193.400 36.755 194.540 ;
        RECT 36.925 193.570 37.255 194.550 ;
        RECT 37.425 193.400 37.635 194.540 ;
        RECT 37.865 194.370 38.135 195.380 ;
        RECT 38.305 195.210 39.530 195.380 ;
        RECT 39.705 195.225 39.995 195.950 ;
        RECT 40.170 195.320 40.505 195.780 ;
        RECT 40.675 195.490 40.845 195.950 ;
        RECT 41.015 195.320 41.345 195.780 ;
        RECT 41.515 195.490 41.685 195.950 ;
        RECT 41.855 195.570 43.865 195.780 ;
        RECT 41.855 195.320 42.105 195.570 ;
        RECT 38.305 194.540 38.475 195.210 ;
        RECT 40.170 195.130 42.105 195.320 ;
        RECT 42.275 195.230 43.445 195.400 ;
        RECT 38.645 194.710 39.025 195.040 ;
        RECT 39.195 194.710 39.530 195.040 ;
        RECT 42.275 194.960 42.525 195.230 ;
        RECT 43.615 195.150 43.865 195.570 ;
        RECT 44.320 195.380 44.575 195.730 ;
        RECT 44.745 195.550 45.075 195.950 ;
        RECT 45.245 195.380 45.415 195.730 ;
        RECT 45.585 195.550 45.965 195.950 ;
        RECT 44.320 195.210 45.985 195.380 ;
        RECT 46.155 195.275 46.430 195.620 ;
        RECT 45.815 195.040 45.985 195.210 ;
        RECT 40.190 194.710 41.810 194.960 ;
        RECT 38.305 194.370 38.620 194.540 ;
        RECT 37.870 193.400 38.185 194.200 ;
        RECT 38.450 193.755 38.620 194.370 ;
        RECT 38.790 194.030 39.025 194.710 ;
        RECT 39.195 193.755 39.530 194.540 ;
        RECT 38.450 193.585 39.530 193.755 ;
        RECT 39.705 193.400 39.995 194.565 ;
        RECT 41.990 194.540 42.525 194.960 ;
        RECT 42.695 194.710 44.135 194.960 ;
        RECT 44.305 194.710 44.650 195.040 ;
        RECT 44.820 194.710 45.645 195.040 ;
        RECT 45.815 194.710 46.090 195.040 ;
        RECT 40.170 193.400 40.425 194.540 ;
        RECT 40.595 194.370 43.445 194.540 ;
        RECT 40.595 193.570 40.925 194.370 ;
        RECT 41.095 193.400 41.265 194.200 ;
        RECT 41.435 193.570 41.765 194.370 ;
        RECT 41.935 193.400 42.105 194.200 ;
        RECT 42.275 193.570 42.605 194.370 ;
        RECT 42.775 193.400 42.945 194.200 ;
        RECT 43.115 193.570 43.445 194.370 ;
        RECT 44.325 194.250 44.650 194.540 ;
        RECT 44.820 194.420 45.015 194.710 ;
        RECT 45.815 194.540 45.985 194.710 ;
        RECT 46.260 194.540 46.430 195.275 ;
        RECT 46.605 195.150 47.300 195.780 ;
        RECT 47.505 195.150 47.815 195.950 ;
        RECT 46.625 194.710 46.960 194.960 ;
        RECT 47.130 194.550 47.300 195.150 ;
        RECT 48.260 195.140 48.505 195.745 ;
        RECT 48.725 195.415 49.235 195.950 ;
        RECT 47.470 194.710 47.805 194.980 ;
        RECT 47.985 194.970 49.215 195.140 ;
        RECT 45.325 194.370 45.985 194.540 ;
        RECT 45.325 194.250 45.495 194.370 ;
        RECT 43.615 193.400 43.865 194.200 ;
        RECT 44.325 194.080 45.495 194.250 ;
        RECT 44.305 193.620 45.495 193.910 ;
        RECT 45.665 193.400 45.945 194.200 ;
        RECT 46.155 193.570 46.430 194.540 ;
        RECT 46.605 193.400 46.865 194.540 ;
        RECT 47.035 193.570 47.365 194.550 ;
        RECT 47.535 193.400 47.815 194.540 ;
        RECT 47.985 194.160 48.325 194.970 ;
        RECT 48.495 194.405 49.245 194.595 ;
        RECT 47.985 193.750 48.500 194.160 ;
        RECT 48.735 193.400 48.905 194.160 ;
        RECT 49.075 193.740 49.245 194.405 ;
        RECT 49.415 194.420 49.605 195.780 ;
        RECT 49.775 195.610 50.050 195.780 ;
        RECT 49.775 195.440 50.055 195.610 ;
        RECT 49.775 194.620 50.050 195.440 ;
        RECT 50.240 195.415 50.770 195.780 ;
        RECT 51.195 195.550 51.525 195.950 ;
        RECT 50.595 195.380 50.770 195.415 ;
        RECT 50.255 194.420 50.425 195.220 ;
        RECT 49.415 194.250 50.425 194.420 ;
        RECT 50.595 195.210 51.525 195.380 ;
        RECT 51.695 195.210 51.950 195.780 ;
        RECT 50.595 194.080 50.765 195.210 ;
        RECT 51.355 195.040 51.525 195.210 ;
        RECT 49.640 193.910 50.765 194.080 ;
        RECT 50.935 194.710 51.130 195.040 ;
        RECT 51.355 194.710 51.610 195.040 ;
        RECT 50.935 193.740 51.105 194.710 ;
        RECT 51.780 194.540 51.950 195.210 ;
        RECT 49.075 193.570 51.105 193.740 ;
        RECT 51.275 193.400 51.445 194.540 ;
        RECT 51.615 193.570 51.950 194.540 ;
        RECT 52.135 195.225 52.465 195.735 ;
        RECT 52.635 195.550 52.965 195.950 ;
        RECT 54.015 195.380 54.345 195.720 ;
        RECT 54.515 195.550 54.845 195.950 ;
        RECT 52.135 194.460 52.325 195.225 ;
        RECT 52.635 195.210 55.000 195.380 ;
        RECT 52.635 195.040 52.805 195.210 ;
        RECT 52.495 194.710 52.805 195.040 ;
        RECT 52.975 194.710 53.280 195.040 ;
        RECT 52.135 193.610 52.465 194.460 ;
        RECT 52.635 193.400 52.885 194.540 ;
        RECT 53.065 194.380 53.280 194.710 ;
        RECT 53.455 194.380 53.740 195.040 ;
        RECT 53.935 194.380 54.200 195.040 ;
        RECT 54.415 194.380 54.660 195.040 ;
        RECT 54.830 194.210 55.000 195.210 ;
        RECT 55.350 195.185 55.805 195.950 ;
        RECT 56.080 195.570 57.380 195.780 ;
        RECT 57.635 195.590 57.965 195.950 ;
        RECT 57.210 195.420 57.380 195.570 ;
        RECT 58.135 195.450 58.395 195.780 ;
        RECT 56.280 194.960 56.500 195.360 ;
        RECT 55.345 194.760 55.835 194.960 ;
        RECT 56.025 194.750 56.500 194.960 ;
        RECT 56.745 194.960 56.955 195.360 ;
        RECT 57.210 195.295 57.965 195.420 ;
        RECT 57.210 195.250 58.055 195.295 ;
        RECT 57.785 195.130 58.055 195.250 ;
        RECT 56.745 194.750 57.075 194.960 ;
        RECT 57.245 194.690 57.655 194.995 ;
        RECT 53.075 194.040 54.365 194.210 ;
        RECT 53.075 193.620 53.325 194.040 ;
        RECT 53.555 193.400 53.885 193.870 ;
        RECT 54.115 193.620 54.365 194.040 ;
        RECT 54.545 194.040 55.000 194.210 ;
        RECT 55.350 194.520 56.525 194.580 ;
        RECT 57.885 194.555 58.055 195.130 ;
        RECT 57.855 194.520 58.055 194.555 ;
        RECT 55.350 194.410 58.055 194.520 ;
        RECT 54.545 193.610 54.875 194.040 ;
        RECT 55.350 193.790 55.605 194.410 ;
        RECT 56.195 194.350 57.995 194.410 ;
        RECT 56.195 194.320 56.525 194.350 ;
        RECT 58.225 194.250 58.395 195.450 ;
        RECT 58.570 195.185 59.025 195.950 ;
        RECT 59.300 195.570 60.600 195.780 ;
        RECT 60.855 195.590 61.185 195.950 ;
        RECT 60.430 195.420 60.600 195.570 ;
        RECT 61.355 195.450 61.615 195.780 ;
        RECT 61.385 195.440 61.615 195.450 ;
        RECT 59.500 194.960 59.720 195.360 ;
        RECT 58.565 194.760 59.055 194.960 ;
        RECT 59.245 194.750 59.720 194.960 ;
        RECT 59.965 194.960 60.175 195.360 ;
        RECT 60.430 195.295 61.185 195.420 ;
        RECT 60.430 195.250 61.275 195.295 ;
        RECT 61.005 195.130 61.275 195.250 ;
        RECT 59.965 194.750 60.295 194.960 ;
        RECT 60.465 194.690 60.875 194.995 ;
        RECT 55.855 194.150 56.040 194.240 ;
        RECT 56.630 194.150 57.465 194.160 ;
        RECT 55.855 193.950 57.465 194.150 ;
        RECT 55.855 193.910 56.085 193.950 ;
        RECT 55.350 193.570 55.685 193.790 ;
        RECT 56.690 193.400 57.045 193.780 ;
        RECT 57.215 193.570 57.465 193.950 ;
        RECT 57.715 193.400 57.965 194.180 ;
        RECT 58.135 193.570 58.395 194.250 ;
        RECT 58.570 194.520 59.745 194.580 ;
        RECT 61.105 194.555 61.275 195.130 ;
        RECT 61.075 194.520 61.275 194.555 ;
        RECT 58.570 194.410 61.275 194.520 ;
        RECT 58.570 193.790 58.825 194.410 ;
        RECT 59.415 194.350 61.215 194.410 ;
        RECT 59.415 194.320 59.745 194.350 ;
        RECT 61.445 194.250 61.615 195.440 ;
        RECT 61.785 195.180 65.295 195.950 ;
        RECT 65.465 195.225 65.755 195.950 ;
        RECT 65.930 195.185 66.385 195.950 ;
        RECT 66.660 195.570 67.960 195.780 ;
        RECT 68.215 195.590 68.545 195.950 ;
        RECT 67.790 195.420 67.960 195.570 ;
        RECT 68.715 195.450 68.975 195.780 ;
        RECT 61.785 194.660 63.435 195.180 ;
        RECT 63.605 194.490 65.295 195.010 ;
        RECT 66.860 194.960 67.080 195.360 ;
        RECT 65.925 194.760 66.415 194.960 ;
        RECT 66.605 194.750 67.080 194.960 ;
        RECT 67.325 194.960 67.535 195.360 ;
        RECT 67.790 195.295 68.545 195.420 ;
        RECT 67.790 195.250 68.635 195.295 ;
        RECT 68.365 195.130 68.635 195.250 ;
        RECT 67.325 194.750 67.655 194.960 ;
        RECT 67.825 194.690 68.235 194.995 ;
        RECT 59.075 194.150 59.260 194.240 ;
        RECT 59.850 194.150 60.685 194.160 ;
        RECT 59.075 193.950 60.685 194.150 ;
        RECT 59.075 193.910 59.305 193.950 ;
        RECT 58.570 193.570 58.905 193.790 ;
        RECT 59.910 193.400 60.265 193.780 ;
        RECT 60.435 193.570 60.685 193.950 ;
        RECT 60.935 193.400 61.185 194.180 ;
        RECT 61.355 193.570 61.615 194.250 ;
        RECT 61.785 193.400 65.295 194.490 ;
        RECT 65.465 193.400 65.755 194.565 ;
        RECT 65.930 194.520 67.105 194.580 ;
        RECT 68.465 194.555 68.635 195.130 ;
        RECT 68.435 194.520 68.635 194.555 ;
        RECT 65.930 194.410 68.635 194.520 ;
        RECT 65.930 193.790 66.185 194.410 ;
        RECT 66.775 194.350 68.575 194.410 ;
        RECT 66.775 194.320 67.105 194.350 ;
        RECT 68.805 194.250 68.975 195.450 ;
        RECT 69.150 195.400 69.405 195.690 ;
        RECT 69.575 195.570 69.905 195.950 ;
        RECT 69.150 195.230 69.900 195.400 ;
        RECT 69.150 194.410 69.500 195.060 ;
        RECT 66.435 194.150 66.620 194.240 ;
        RECT 67.210 194.150 68.045 194.160 ;
        RECT 66.435 193.950 68.045 194.150 ;
        RECT 66.435 193.910 66.665 193.950 ;
        RECT 65.930 193.570 66.265 193.790 ;
        RECT 67.270 193.400 67.625 193.780 ;
        RECT 67.795 193.570 68.045 193.950 ;
        RECT 68.295 193.400 68.545 194.180 ;
        RECT 68.715 193.570 68.975 194.250 ;
        RECT 69.670 194.240 69.900 195.230 ;
        RECT 69.150 194.070 69.900 194.240 ;
        RECT 69.150 193.570 69.405 194.070 ;
        RECT 69.575 193.400 69.905 193.900 ;
        RECT 70.075 193.570 70.245 195.690 ;
        RECT 70.605 195.590 70.935 195.950 ;
        RECT 71.105 195.560 71.600 195.730 ;
        RECT 71.805 195.560 72.660 195.730 ;
        RECT 70.475 194.370 70.935 195.420 ;
        RECT 70.415 193.585 70.740 194.370 ;
        RECT 71.105 194.200 71.275 195.560 ;
        RECT 71.445 194.650 71.795 195.270 ;
        RECT 71.965 195.050 72.320 195.270 ;
        RECT 71.965 194.460 72.135 195.050 ;
        RECT 72.490 194.850 72.660 195.560 ;
        RECT 73.535 195.490 73.865 195.950 ;
        RECT 74.075 195.590 74.425 195.760 ;
        RECT 72.865 195.020 73.655 195.270 ;
        RECT 74.075 195.200 74.335 195.590 ;
        RECT 74.645 195.500 75.595 195.780 ;
        RECT 75.765 195.510 75.955 195.950 ;
        RECT 76.125 195.570 77.195 195.740 ;
        RECT 73.825 194.850 73.995 195.030 ;
        RECT 71.105 194.030 71.500 194.200 ;
        RECT 71.670 194.070 72.135 194.460 ;
        RECT 72.305 194.680 73.995 194.850 ;
        RECT 71.330 193.900 71.500 194.030 ;
        RECT 72.305 193.900 72.475 194.680 ;
        RECT 74.165 194.510 74.335 195.200 ;
        RECT 72.835 194.340 74.335 194.510 ;
        RECT 74.525 194.540 74.735 195.330 ;
        RECT 74.905 194.710 75.255 195.330 ;
        RECT 75.425 194.720 75.595 195.500 ;
        RECT 76.125 195.340 76.295 195.570 ;
        RECT 75.765 195.170 76.295 195.340 ;
        RECT 75.765 194.890 75.985 195.170 ;
        RECT 76.465 195.000 76.705 195.400 ;
        RECT 75.425 194.550 75.830 194.720 ;
        RECT 76.165 194.630 76.705 195.000 ;
        RECT 76.875 195.215 77.195 195.570 ;
        RECT 76.875 194.960 77.200 195.215 ;
        RECT 77.395 195.140 77.565 195.950 ;
        RECT 77.735 195.300 78.065 195.780 ;
        RECT 78.235 195.480 78.405 195.950 ;
        RECT 78.575 195.300 78.905 195.780 ;
        RECT 79.075 195.480 79.245 195.950 ;
        RECT 80.035 195.480 80.205 195.950 ;
        RECT 80.375 195.300 80.705 195.780 ;
        RECT 80.875 195.480 81.045 195.950 ;
        RECT 81.215 195.300 81.545 195.780 ;
        RECT 77.735 195.130 79.500 195.300 ;
        RECT 76.875 194.750 78.905 194.960 ;
        RECT 76.875 194.740 77.220 194.750 ;
        RECT 74.525 194.380 75.200 194.540 ;
        RECT 75.660 194.460 75.830 194.550 ;
        RECT 74.525 194.370 75.490 194.380 ;
        RECT 74.165 194.200 74.335 194.340 ;
        RECT 70.910 193.400 71.160 193.860 ;
        RECT 71.330 193.570 71.580 193.900 ;
        RECT 71.795 193.570 72.475 193.900 ;
        RECT 72.645 194.000 73.720 194.170 ;
        RECT 74.165 194.030 74.725 194.200 ;
        RECT 75.030 194.080 75.490 194.370 ;
        RECT 75.660 194.290 76.880 194.460 ;
        RECT 72.645 193.660 72.815 194.000 ;
        RECT 73.050 193.400 73.380 193.830 ;
        RECT 73.550 193.660 73.720 194.000 ;
        RECT 74.015 193.400 74.385 193.860 ;
        RECT 74.555 193.570 74.725 194.030 ;
        RECT 75.660 193.910 75.830 194.290 ;
        RECT 77.050 194.120 77.220 194.740 ;
        RECT 79.090 194.580 79.500 195.130 ;
        RECT 74.960 193.570 75.830 193.910 ;
        RECT 76.420 193.950 77.220 194.120 ;
        RECT 76.000 193.400 76.250 193.860 ;
        RECT 76.420 193.660 76.590 193.950 ;
        RECT 76.770 193.400 77.100 193.780 ;
        RECT 77.395 193.400 77.565 194.460 ;
        RECT 77.775 194.410 79.500 194.580 ;
        RECT 79.780 195.130 81.545 195.300 ;
        RECT 81.715 195.140 81.885 195.950 ;
        RECT 82.085 195.570 83.155 195.740 ;
        RECT 82.085 195.215 82.405 195.570 ;
        RECT 79.780 194.580 80.190 195.130 ;
        RECT 82.080 194.960 82.405 195.215 ;
        RECT 80.375 194.750 82.405 194.960 ;
        RECT 82.060 194.740 82.405 194.750 ;
        RECT 82.575 195.000 82.815 195.400 ;
        RECT 82.985 195.340 83.155 195.570 ;
        RECT 83.325 195.510 83.515 195.950 ;
        RECT 83.685 195.500 84.635 195.780 ;
        RECT 84.855 195.590 85.205 195.760 ;
        RECT 82.985 195.170 83.515 195.340 ;
        RECT 79.780 194.410 81.505 194.580 ;
        RECT 77.775 193.570 78.065 194.410 ;
        RECT 78.235 193.400 78.405 194.240 ;
        RECT 78.615 193.570 78.865 194.410 ;
        RECT 79.075 193.400 79.245 194.240 ;
        RECT 80.035 193.400 80.205 194.240 ;
        RECT 80.415 193.570 80.665 194.410 ;
        RECT 80.875 193.400 81.045 194.240 ;
        RECT 81.215 193.570 81.505 194.410 ;
        RECT 81.715 193.400 81.885 194.460 ;
        RECT 82.060 194.120 82.230 194.740 ;
        RECT 82.575 194.630 83.115 195.000 ;
        RECT 83.295 194.890 83.515 195.170 ;
        RECT 83.685 194.720 83.855 195.500 ;
        RECT 83.450 194.550 83.855 194.720 ;
        RECT 84.025 194.710 84.375 195.330 ;
        RECT 83.450 194.460 83.620 194.550 ;
        RECT 84.545 194.540 84.755 195.330 ;
        RECT 82.400 194.290 83.620 194.460 ;
        RECT 84.080 194.380 84.755 194.540 ;
        RECT 82.060 193.950 82.860 194.120 ;
        RECT 82.180 193.400 82.510 193.780 ;
        RECT 82.690 193.660 82.860 193.950 ;
        RECT 83.450 193.910 83.620 194.290 ;
        RECT 83.790 194.370 84.755 194.380 ;
        RECT 84.945 195.200 85.205 195.590 ;
        RECT 85.415 195.490 85.745 195.950 ;
        RECT 86.620 195.560 87.475 195.730 ;
        RECT 87.680 195.560 88.175 195.730 ;
        RECT 88.345 195.590 88.675 195.950 ;
        RECT 84.945 194.510 85.115 195.200 ;
        RECT 85.285 194.850 85.455 195.030 ;
        RECT 85.625 195.020 86.415 195.270 ;
        RECT 86.620 194.850 86.790 195.560 ;
        RECT 86.960 195.050 87.315 195.270 ;
        RECT 85.285 194.680 86.975 194.850 ;
        RECT 83.790 194.080 84.250 194.370 ;
        RECT 84.945 194.340 86.445 194.510 ;
        RECT 84.945 194.200 85.115 194.340 ;
        RECT 84.555 194.030 85.115 194.200 ;
        RECT 83.030 193.400 83.280 193.860 ;
        RECT 83.450 193.570 84.320 193.910 ;
        RECT 84.555 193.570 84.725 194.030 ;
        RECT 85.560 194.000 86.635 194.170 ;
        RECT 84.895 193.400 85.265 193.860 ;
        RECT 85.560 193.660 85.730 194.000 ;
        RECT 85.900 193.400 86.230 193.830 ;
        RECT 86.465 193.660 86.635 194.000 ;
        RECT 86.805 193.900 86.975 194.680 ;
        RECT 87.145 194.460 87.315 195.050 ;
        RECT 87.485 194.650 87.835 195.270 ;
        RECT 87.145 194.070 87.610 194.460 ;
        RECT 88.005 194.200 88.175 195.560 ;
        RECT 88.345 194.370 88.805 195.420 ;
        RECT 87.780 194.030 88.175 194.200 ;
        RECT 87.780 193.900 87.950 194.030 ;
        RECT 86.805 193.570 87.485 193.900 ;
        RECT 87.700 193.570 87.950 193.900 ;
        RECT 88.120 193.400 88.370 193.860 ;
        RECT 88.540 193.585 88.865 194.370 ;
        RECT 89.035 193.570 89.205 195.690 ;
        RECT 89.375 195.570 89.705 195.950 ;
        RECT 89.875 195.400 90.130 195.690 ;
        RECT 89.380 195.230 90.130 195.400 ;
        RECT 89.380 194.240 89.610 195.230 ;
        RECT 91.225 195.225 91.515 195.950 ;
        RECT 91.690 195.400 91.945 195.690 ;
        RECT 92.115 195.570 92.445 195.950 ;
        RECT 91.690 195.230 92.440 195.400 ;
        RECT 89.780 194.410 90.130 195.060 ;
        RECT 89.380 194.070 90.130 194.240 ;
        RECT 89.375 193.400 89.705 193.900 ;
        RECT 89.875 193.570 90.130 194.070 ;
        RECT 91.225 193.400 91.515 194.565 ;
        RECT 91.690 194.410 92.040 195.060 ;
        RECT 92.210 194.240 92.440 195.230 ;
        RECT 91.690 194.070 92.440 194.240 ;
        RECT 91.690 193.570 91.945 194.070 ;
        RECT 92.115 193.400 92.445 193.900 ;
        RECT 92.615 193.570 92.785 195.690 ;
        RECT 93.145 195.590 93.475 195.950 ;
        RECT 93.645 195.560 94.140 195.730 ;
        RECT 94.345 195.560 95.200 195.730 ;
        RECT 93.015 194.370 93.475 195.420 ;
        RECT 92.955 193.585 93.280 194.370 ;
        RECT 93.645 194.200 93.815 195.560 ;
        RECT 93.985 194.650 94.335 195.270 ;
        RECT 94.505 195.050 94.860 195.270 ;
        RECT 94.505 194.460 94.675 195.050 ;
        RECT 95.030 194.850 95.200 195.560 ;
        RECT 96.075 195.490 96.405 195.950 ;
        RECT 96.615 195.590 96.965 195.760 ;
        RECT 95.405 195.020 96.195 195.270 ;
        RECT 96.615 195.200 96.875 195.590 ;
        RECT 97.185 195.500 98.135 195.780 ;
        RECT 98.305 195.510 98.495 195.950 ;
        RECT 98.665 195.570 99.735 195.740 ;
        RECT 96.365 194.850 96.535 195.030 ;
        RECT 93.645 194.030 94.040 194.200 ;
        RECT 94.210 194.070 94.675 194.460 ;
        RECT 94.845 194.680 96.535 194.850 ;
        RECT 93.870 193.900 94.040 194.030 ;
        RECT 94.845 193.900 95.015 194.680 ;
        RECT 96.705 194.510 96.875 195.200 ;
        RECT 95.375 194.340 96.875 194.510 ;
        RECT 97.065 194.540 97.275 195.330 ;
        RECT 97.445 194.710 97.795 195.330 ;
        RECT 97.965 194.720 98.135 195.500 ;
        RECT 98.665 195.340 98.835 195.570 ;
        RECT 98.305 195.170 98.835 195.340 ;
        RECT 98.305 194.890 98.525 195.170 ;
        RECT 99.005 195.000 99.245 195.400 ;
        RECT 97.965 194.550 98.370 194.720 ;
        RECT 98.705 194.630 99.245 195.000 ;
        RECT 99.415 195.215 99.735 195.570 ;
        RECT 99.415 194.960 99.740 195.215 ;
        RECT 99.935 195.140 100.105 195.950 ;
        RECT 100.275 195.300 100.605 195.780 ;
        RECT 100.775 195.480 100.945 195.950 ;
        RECT 101.115 195.300 101.445 195.780 ;
        RECT 101.615 195.480 101.785 195.950 ;
        RECT 100.275 195.130 102.040 195.300 ;
        RECT 99.415 194.750 101.445 194.960 ;
        RECT 99.415 194.740 99.760 194.750 ;
        RECT 97.065 194.380 97.740 194.540 ;
        RECT 98.200 194.460 98.370 194.550 ;
        RECT 97.065 194.370 98.030 194.380 ;
        RECT 96.705 194.200 96.875 194.340 ;
        RECT 93.450 193.400 93.700 193.860 ;
        RECT 93.870 193.570 94.120 193.900 ;
        RECT 94.335 193.570 95.015 193.900 ;
        RECT 95.185 194.000 96.260 194.170 ;
        RECT 96.705 194.030 97.265 194.200 ;
        RECT 97.570 194.080 98.030 194.370 ;
        RECT 98.200 194.290 99.420 194.460 ;
        RECT 95.185 193.660 95.355 194.000 ;
        RECT 95.590 193.400 95.920 193.830 ;
        RECT 96.090 193.660 96.260 194.000 ;
        RECT 96.555 193.400 96.925 193.860 ;
        RECT 97.095 193.570 97.265 194.030 ;
        RECT 98.200 193.910 98.370 194.290 ;
        RECT 99.590 194.120 99.760 194.740 ;
        RECT 101.630 194.580 102.040 195.130 ;
        RECT 97.500 193.570 98.370 193.910 ;
        RECT 98.960 193.950 99.760 194.120 ;
        RECT 98.540 193.400 98.790 193.860 ;
        RECT 98.960 193.660 99.130 193.950 ;
        RECT 99.310 193.400 99.640 193.780 ;
        RECT 99.935 193.400 100.105 194.460 ;
        RECT 100.315 194.410 102.040 194.580 ;
        RECT 102.265 195.275 102.525 195.780 ;
        RECT 102.705 195.570 103.035 195.950 ;
        RECT 103.215 195.400 103.385 195.780 ;
        RECT 102.265 194.475 102.435 195.275 ;
        RECT 102.720 195.230 103.385 195.400 ;
        RECT 102.720 194.975 102.890 195.230 ;
        RECT 103.665 195.140 103.905 195.950 ;
        RECT 104.075 195.140 104.405 195.780 ;
        RECT 104.575 195.140 104.845 195.950 ;
        RECT 105.945 195.275 106.205 195.780 ;
        RECT 106.385 195.570 106.715 195.950 ;
        RECT 106.895 195.400 107.065 195.780 ;
        RECT 102.605 194.645 102.890 194.975 ;
        RECT 103.125 194.680 103.455 195.050 ;
        RECT 103.645 194.710 103.995 194.960 ;
        RECT 102.720 194.500 102.890 194.645 ;
        RECT 104.165 194.540 104.335 195.140 ;
        RECT 104.505 194.710 104.855 194.960 ;
        RECT 100.315 193.570 100.605 194.410 ;
        RECT 100.775 193.400 100.945 194.240 ;
        RECT 101.155 193.570 101.405 194.410 ;
        RECT 101.615 193.400 101.785 194.240 ;
        RECT 102.265 193.570 102.535 194.475 ;
        RECT 102.720 194.330 103.385 194.500 ;
        RECT 102.705 193.400 103.035 194.160 ;
        RECT 103.215 193.570 103.385 194.330 ;
        RECT 103.655 194.370 104.335 194.540 ;
        RECT 103.655 193.585 103.985 194.370 ;
        RECT 104.515 193.400 104.845 194.540 ;
        RECT 105.945 194.475 106.115 195.275 ;
        RECT 106.400 195.230 107.065 195.400 ;
        RECT 106.400 194.975 106.570 195.230 ;
        RECT 107.325 195.115 107.615 195.950 ;
        RECT 107.785 195.550 108.740 195.720 ;
        RECT 109.155 195.560 109.485 195.950 ;
        RECT 106.285 194.645 106.570 194.975 ;
        RECT 106.805 194.680 107.135 195.050 ;
        RECT 107.785 194.670 107.955 195.550 ;
        RECT 109.655 195.380 109.825 195.700 ;
        RECT 109.995 195.560 110.325 195.950 ;
        RECT 108.125 195.210 110.375 195.380 ;
        RECT 111.025 195.220 111.315 195.950 ;
        RECT 108.125 194.710 108.355 195.210 ;
        RECT 108.525 194.790 108.900 194.960 ;
        RECT 106.400 194.500 106.570 194.645 ;
        RECT 107.325 194.500 107.955 194.670 ;
        RECT 108.730 194.590 108.900 194.790 ;
        RECT 109.070 194.760 109.620 194.960 ;
        RECT 109.790 194.590 110.035 195.040 ;
        RECT 105.945 193.570 106.215 194.475 ;
        RECT 106.400 194.330 107.065 194.500 ;
        RECT 106.385 193.400 106.715 194.160 ;
        RECT 106.895 193.570 107.065 194.330 ;
        RECT 107.325 193.570 107.645 194.500 ;
        RECT 108.730 194.420 110.035 194.590 ;
        RECT 110.205 194.250 110.375 195.210 ;
        RECT 111.015 194.710 111.315 195.040 ;
        RECT 111.495 195.020 111.725 195.660 ;
        RECT 111.905 195.400 112.215 195.770 ;
        RECT 112.395 195.580 113.065 195.950 ;
        RECT 111.905 195.200 113.135 195.400 ;
        RECT 111.495 194.710 112.020 195.020 ;
        RECT 112.200 194.710 112.665 195.020 ;
        RECT 112.845 194.530 113.135 195.200 ;
        RECT 107.825 194.080 109.065 194.250 ;
        RECT 107.825 193.570 108.225 194.080 ;
        RECT 108.395 193.400 108.565 193.910 ;
        RECT 108.735 193.570 109.065 194.080 ;
        RECT 109.235 193.400 109.405 194.250 ;
        RECT 109.995 193.570 110.375 194.250 ;
        RECT 111.025 194.290 112.185 194.530 ;
        RECT 111.025 193.580 111.285 194.290 ;
        RECT 111.455 193.400 111.785 194.110 ;
        RECT 111.955 193.580 112.185 194.290 ;
        RECT 112.365 194.310 113.135 194.530 ;
        RECT 112.365 193.580 112.635 194.310 ;
        RECT 112.815 193.400 113.155 194.130 ;
        RECT 113.325 193.580 113.585 195.770 ;
        RECT 113.770 195.185 114.225 195.950 ;
        RECT 114.500 195.570 115.800 195.780 ;
        RECT 116.055 195.590 116.385 195.950 ;
        RECT 115.630 195.420 115.800 195.570 ;
        RECT 116.555 195.450 116.815 195.780 ;
        RECT 114.700 194.960 114.920 195.360 ;
        RECT 113.765 194.760 114.255 194.960 ;
        RECT 114.445 194.750 114.920 194.960 ;
        RECT 115.165 194.960 115.375 195.360 ;
        RECT 115.630 195.295 116.385 195.420 ;
        RECT 115.630 195.250 116.475 195.295 ;
        RECT 116.205 195.130 116.475 195.250 ;
        RECT 115.165 194.750 115.495 194.960 ;
        RECT 115.665 194.690 116.075 194.995 ;
        RECT 113.770 194.520 114.945 194.580 ;
        RECT 116.305 194.555 116.475 195.130 ;
        RECT 116.275 194.520 116.475 194.555 ;
        RECT 113.770 194.410 116.475 194.520 ;
        RECT 113.770 193.790 114.025 194.410 ;
        RECT 114.615 194.350 116.415 194.410 ;
        RECT 114.615 194.320 114.945 194.350 ;
        RECT 116.645 194.250 116.815 195.450 ;
        RECT 116.985 195.225 117.275 195.950 ;
        RECT 117.445 195.380 117.965 195.780 ;
        RECT 118.135 195.550 118.465 195.950 ;
        RECT 118.635 195.380 118.805 195.725 ;
        RECT 117.445 195.210 118.805 195.380 ;
        RECT 118.975 195.210 119.305 195.950 ;
        RECT 119.540 195.380 119.710 195.630 ;
        RECT 120.210 195.400 120.465 195.690 ;
        RECT 120.635 195.570 120.965 195.950 ;
        RECT 119.540 195.210 120.035 195.380 ;
        RECT 120.210 195.230 120.960 195.400 ;
        RECT 117.445 194.590 117.615 195.210 ;
        RECT 117.785 194.790 118.245 194.960 ;
        RECT 114.275 194.150 114.460 194.240 ;
        RECT 115.050 194.150 115.885 194.160 ;
        RECT 114.275 193.950 115.885 194.150 ;
        RECT 114.275 193.910 114.505 193.950 ;
        RECT 113.770 193.570 114.105 193.790 ;
        RECT 115.110 193.400 115.465 193.780 ;
        RECT 115.635 193.570 115.885 193.950 ;
        RECT 116.135 193.400 116.385 194.180 ;
        RECT 116.555 193.570 116.815 194.250 ;
        RECT 116.985 193.400 117.275 194.565 ;
        RECT 117.445 193.580 117.905 194.590 ;
        RECT 118.075 194.250 118.245 194.790 ;
        RECT 118.425 194.420 118.665 195.040 ;
        RECT 118.835 194.420 119.175 195.040 ;
        RECT 119.345 194.420 119.695 195.040 ;
        RECT 119.865 194.250 120.035 195.210 ;
        RECT 120.210 194.410 120.560 195.060 ;
        RECT 118.075 194.080 120.035 194.250 ;
        RECT 120.730 194.240 120.960 195.230 ;
        RECT 120.210 194.070 120.960 194.240 ;
        RECT 118.975 193.400 119.305 193.910 ;
        RECT 120.210 193.570 120.465 194.070 ;
        RECT 120.635 193.400 120.965 193.900 ;
        RECT 121.135 193.570 121.305 195.690 ;
        RECT 121.665 195.590 121.995 195.950 ;
        RECT 122.165 195.560 122.660 195.730 ;
        RECT 122.865 195.560 123.720 195.730 ;
        RECT 121.535 194.370 121.995 195.420 ;
        RECT 121.475 193.585 121.800 194.370 ;
        RECT 122.165 194.200 122.335 195.560 ;
        RECT 122.505 194.650 122.855 195.270 ;
        RECT 123.025 195.050 123.380 195.270 ;
        RECT 123.025 194.460 123.195 195.050 ;
        RECT 123.550 194.850 123.720 195.560 ;
        RECT 124.595 195.490 124.925 195.950 ;
        RECT 125.135 195.590 125.485 195.760 ;
        RECT 123.925 195.020 124.715 195.270 ;
        RECT 125.135 195.200 125.395 195.590 ;
        RECT 125.705 195.500 126.655 195.780 ;
        RECT 126.825 195.510 127.015 195.950 ;
        RECT 127.185 195.570 128.255 195.740 ;
        RECT 124.885 194.850 125.055 195.030 ;
        RECT 122.165 194.030 122.560 194.200 ;
        RECT 122.730 194.070 123.195 194.460 ;
        RECT 123.365 194.680 125.055 194.850 ;
        RECT 122.390 193.900 122.560 194.030 ;
        RECT 123.365 193.900 123.535 194.680 ;
        RECT 125.225 194.510 125.395 195.200 ;
        RECT 123.895 194.340 125.395 194.510 ;
        RECT 125.585 194.540 125.795 195.330 ;
        RECT 125.965 194.710 126.315 195.330 ;
        RECT 126.485 194.720 126.655 195.500 ;
        RECT 127.185 195.340 127.355 195.570 ;
        RECT 126.825 195.170 127.355 195.340 ;
        RECT 126.825 194.890 127.045 195.170 ;
        RECT 127.525 195.000 127.765 195.400 ;
        RECT 126.485 194.550 126.890 194.720 ;
        RECT 127.225 194.630 127.765 195.000 ;
        RECT 127.935 195.215 128.255 195.570 ;
        RECT 128.500 195.490 128.805 195.950 ;
        RECT 128.975 195.240 129.230 195.770 ;
        RECT 127.935 195.040 128.260 195.215 ;
        RECT 127.935 194.740 128.850 195.040 ;
        RECT 128.110 194.710 128.850 194.740 ;
        RECT 125.585 194.380 126.260 194.540 ;
        RECT 126.720 194.460 126.890 194.550 ;
        RECT 125.585 194.370 126.550 194.380 ;
        RECT 125.225 194.200 125.395 194.340 ;
        RECT 121.970 193.400 122.220 193.860 ;
        RECT 122.390 193.570 122.640 193.900 ;
        RECT 122.855 193.570 123.535 193.900 ;
        RECT 123.705 194.000 124.780 194.170 ;
        RECT 125.225 194.030 125.785 194.200 ;
        RECT 126.090 194.080 126.550 194.370 ;
        RECT 126.720 194.290 127.940 194.460 ;
        RECT 123.705 193.660 123.875 194.000 ;
        RECT 124.110 193.400 124.440 193.830 ;
        RECT 124.610 193.660 124.780 194.000 ;
        RECT 125.075 193.400 125.445 193.860 ;
        RECT 125.615 193.570 125.785 194.030 ;
        RECT 126.720 193.910 126.890 194.290 ;
        RECT 128.110 194.120 128.280 194.710 ;
        RECT 129.020 194.590 129.230 195.240 ;
        RECT 129.405 195.150 129.700 195.950 ;
        RECT 129.870 195.040 130.145 195.780 ;
        RECT 130.315 195.210 130.985 195.950 ;
        RECT 131.155 195.380 131.440 195.725 ;
        RECT 131.620 195.550 131.995 195.950 ;
        RECT 132.210 195.380 132.540 195.725 ;
        RECT 131.155 195.210 132.540 195.380 ;
        RECT 132.790 195.210 133.375 195.780 ;
        RECT 133.565 195.220 133.855 195.950 ;
        RECT 129.870 194.980 130.225 195.040 ;
        RECT 129.405 194.720 130.225 194.980 ;
        RECT 126.020 193.570 126.890 193.910 ;
        RECT 127.480 193.950 128.280 194.120 ;
        RECT 127.060 193.400 127.310 193.860 ;
        RECT 127.480 193.660 127.650 193.950 ;
        RECT 127.830 193.400 128.160 193.780 ;
        RECT 128.500 193.400 128.805 194.540 ;
        RECT 128.975 193.710 129.230 194.590 ;
        RECT 129.405 193.400 129.700 194.550 ;
        RECT 129.870 193.570 130.225 194.720 ;
        RECT 130.395 194.540 130.565 195.040 ;
        RECT 130.735 194.710 131.070 195.040 ;
        RECT 131.240 194.710 131.570 195.040 ;
        RECT 130.395 194.370 131.130 194.540 ;
        RECT 130.395 193.400 130.790 194.200 ;
        RECT 130.960 193.740 131.130 194.370 ;
        RECT 131.300 193.965 131.570 194.710 ;
        RECT 131.760 194.710 132.050 195.040 ;
        RECT 132.220 194.710 132.620 195.040 ;
        RECT 131.760 193.965 131.995 194.710 ;
        RECT 132.790 194.540 132.960 195.210 ;
        RECT 133.130 194.710 133.375 195.040 ;
        RECT 133.555 194.710 133.855 195.040 ;
        RECT 134.035 195.020 134.265 195.660 ;
        RECT 134.445 195.400 134.755 195.770 ;
        RECT 134.935 195.580 135.605 195.950 ;
        RECT 134.445 195.200 135.675 195.400 ;
        RECT 134.035 194.710 134.560 195.020 ;
        RECT 134.740 194.710 135.205 195.020 ;
        RECT 132.165 194.370 133.375 194.540 ;
        RECT 135.385 194.530 135.675 195.200 ;
        RECT 132.165 193.740 132.495 194.370 ;
        RECT 130.960 193.570 132.495 193.740 ;
        RECT 132.680 193.400 132.915 194.200 ;
        RECT 133.085 193.570 133.375 194.370 ;
        RECT 133.565 194.290 134.725 194.530 ;
        RECT 133.565 193.580 133.825 194.290 ;
        RECT 133.995 193.400 134.325 194.110 ;
        RECT 134.495 193.580 134.725 194.290 ;
        RECT 134.905 194.310 135.675 194.530 ;
        RECT 134.905 193.580 135.175 194.310 ;
        RECT 135.355 193.400 135.695 194.130 ;
        RECT 135.865 193.580 136.125 195.770 ;
        RECT 136.310 195.110 136.570 195.950 ;
        RECT 136.745 195.205 137.000 195.780 ;
        RECT 137.170 195.570 137.500 195.950 ;
        RECT 137.715 195.400 137.885 195.780 ;
        RECT 137.170 195.230 137.885 195.400 ;
        RECT 138.235 195.400 138.405 195.780 ;
        RECT 138.620 195.570 138.950 195.950 ;
        RECT 138.235 195.230 138.950 195.400 ;
        RECT 136.310 193.400 136.570 194.550 ;
        RECT 136.745 194.475 136.915 195.205 ;
        RECT 137.170 195.040 137.340 195.230 ;
        RECT 137.085 194.710 137.340 195.040 ;
        RECT 137.170 194.500 137.340 194.710 ;
        RECT 137.620 194.680 137.975 195.050 ;
        RECT 138.145 194.680 138.500 195.050 ;
        RECT 138.780 195.040 138.950 195.230 ;
        RECT 139.120 195.205 139.375 195.780 ;
        RECT 138.780 194.710 139.035 195.040 ;
        RECT 138.780 194.500 138.950 194.710 ;
        RECT 136.745 193.570 137.000 194.475 ;
        RECT 137.170 194.330 137.885 194.500 ;
        RECT 137.170 193.400 137.500 194.160 ;
        RECT 137.715 193.570 137.885 194.330 ;
        RECT 138.235 194.330 138.950 194.500 ;
        RECT 139.205 194.475 139.375 195.205 ;
        RECT 139.550 195.110 139.810 195.950 ;
        RECT 140.995 195.400 141.165 195.780 ;
        RECT 141.380 195.570 141.710 195.950 ;
        RECT 140.995 195.230 141.710 195.400 ;
        RECT 140.905 194.680 141.260 195.050 ;
        RECT 141.540 195.040 141.710 195.230 ;
        RECT 141.880 195.205 142.135 195.780 ;
        RECT 141.540 194.710 141.795 195.040 ;
        RECT 138.235 193.570 138.405 194.330 ;
        RECT 138.620 193.400 138.950 194.160 ;
        RECT 139.120 193.570 139.375 194.475 ;
        RECT 139.550 193.400 139.810 194.550 ;
        RECT 141.540 194.500 141.710 194.710 ;
        RECT 140.995 194.330 141.710 194.500 ;
        RECT 141.965 194.475 142.135 195.205 ;
        RECT 142.310 195.110 142.570 195.950 ;
        RECT 142.745 195.225 143.035 195.950 ;
        RECT 143.225 195.140 143.465 195.950 ;
        RECT 143.635 195.140 143.965 195.780 ;
        RECT 144.135 195.140 144.405 195.950 ;
        RECT 144.675 195.400 144.845 195.780 ;
        RECT 145.060 195.570 145.390 195.950 ;
        RECT 144.675 195.230 145.390 195.400 ;
        RECT 143.205 194.710 143.555 194.960 ;
        RECT 140.995 193.570 141.165 194.330 ;
        RECT 141.380 193.400 141.710 194.160 ;
        RECT 141.880 193.570 142.135 194.475 ;
        RECT 142.310 193.400 142.570 194.550 ;
        RECT 142.745 193.400 143.035 194.565 ;
        RECT 143.725 194.540 143.895 195.140 ;
        RECT 144.065 194.710 144.415 194.960 ;
        RECT 144.585 194.680 144.940 195.050 ;
        RECT 145.220 195.040 145.390 195.230 ;
        RECT 145.560 195.205 145.815 195.780 ;
        RECT 145.220 194.710 145.475 195.040 ;
        RECT 143.215 194.370 143.895 194.540 ;
        RECT 143.215 193.585 143.545 194.370 ;
        RECT 144.075 193.400 144.405 194.540 ;
        RECT 145.220 194.500 145.390 194.710 ;
        RECT 144.675 194.330 145.390 194.500 ;
        RECT 145.645 194.475 145.815 195.205 ;
        RECT 145.990 195.110 146.250 195.950 ;
        RECT 146.425 195.200 147.635 195.950 ;
        RECT 144.675 193.570 144.845 194.330 ;
        RECT 145.060 193.400 145.390 194.160 ;
        RECT 145.560 193.570 145.815 194.475 ;
        RECT 145.990 193.400 146.250 194.550 ;
        RECT 146.425 194.490 146.945 195.030 ;
        RECT 147.115 194.660 147.635 195.200 ;
        RECT 146.425 193.400 147.635 194.490 ;
        RECT 13.860 193.230 147.720 193.400 ;
        RECT 13.945 192.140 15.155 193.230 ;
        RECT 13.945 191.430 14.465 191.970 ;
        RECT 14.635 191.600 15.155 192.140 ;
        RECT 15.330 192.080 15.590 193.230 ;
        RECT 15.765 192.155 16.020 193.060 ;
        RECT 16.190 192.470 16.520 193.230 ;
        RECT 16.735 192.300 16.905 193.060 ;
        RECT 13.945 190.680 15.155 191.430 ;
        RECT 15.330 190.680 15.590 191.520 ;
        RECT 15.765 191.425 15.935 192.155 ;
        RECT 16.190 192.130 16.905 192.300 ;
        RECT 16.190 191.920 16.360 192.130 ;
        RECT 17.170 192.080 17.430 193.230 ;
        RECT 17.605 192.155 17.860 193.060 ;
        RECT 18.030 192.470 18.360 193.230 ;
        RECT 18.575 192.300 18.745 193.060 ;
        RECT 16.105 191.590 16.360 191.920 ;
        RECT 15.765 190.850 16.020 191.425 ;
        RECT 16.190 191.400 16.360 191.590 ;
        RECT 16.640 191.580 16.995 191.950 ;
        RECT 16.190 191.230 16.905 191.400 ;
        RECT 16.190 190.680 16.520 191.060 ;
        RECT 16.735 190.850 16.905 191.230 ;
        RECT 17.170 190.680 17.430 191.520 ;
        RECT 17.605 191.425 17.775 192.155 ;
        RECT 18.030 192.130 18.745 192.300 ;
        RECT 18.030 191.920 18.200 192.130 ;
        RECT 19.010 192.080 19.270 193.230 ;
        RECT 19.445 192.155 19.700 193.060 ;
        RECT 19.870 192.470 20.200 193.230 ;
        RECT 20.415 192.300 20.585 193.060 ;
        RECT 17.945 191.590 18.200 191.920 ;
        RECT 17.605 190.850 17.860 191.425 ;
        RECT 18.030 191.400 18.200 191.590 ;
        RECT 18.480 191.580 18.835 191.950 ;
        RECT 18.030 191.230 18.745 191.400 ;
        RECT 18.030 190.680 18.360 191.060 ;
        RECT 18.575 190.850 18.745 191.230 ;
        RECT 19.010 190.680 19.270 191.520 ;
        RECT 19.445 191.425 19.615 192.155 ;
        RECT 19.870 192.130 20.585 192.300 ;
        RECT 19.870 191.920 20.040 192.130 ;
        RECT 20.850 192.080 21.110 193.230 ;
        RECT 21.285 192.155 21.540 193.060 ;
        RECT 21.710 192.470 22.040 193.230 ;
        RECT 22.255 192.300 22.425 193.060 ;
        RECT 19.785 191.590 20.040 191.920 ;
        RECT 19.445 190.850 19.700 191.425 ;
        RECT 19.870 191.400 20.040 191.590 ;
        RECT 20.320 191.580 20.675 191.950 ;
        RECT 19.870 191.230 20.585 191.400 ;
        RECT 19.870 190.680 20.200 191.060 ;
        RECT 20.415 190.850 20.585 191.230 ;
        RECT 20.850 190.680 21.110 191.520 ;
        RECT 21.285 191.425 21.455 192.155 ;
        RECT 21.710 192.130 22.425 192.300 ;
        RECT 23.145 192.260 23.415 193.030 ;
        RECT 23.585 192.450 23.915 193.230 ;
        RECT 24.120 192.625 24.305 193.030 ;
        RECT 24.475 192.805 24.810 193.230 ;
        RECT 24.120 192.450 24.785 192.625 ;
        RECT 21.710 191.920 21.880 192.130 ;
        RECT 23.145 192.090 24.275 192.260 ;
        RECT 21.625 191.590 21.880 191.920 ;
        RECT 21.285 190.850 21.540 191.425 ;
        RECT 21.710 191.400 21.880 191.590 ;
        RECT 22.160 191.580 22.515 191.950 ;
        RECT 21.710 191.230 22.425 191.400 ;
        RECT 21.710 190.680 22.040 191.060 ;
        RECT 22.255 190.850 22.425 191.230 ;
        RECT 23.145 191.180 23.315 192.090 ;
        RECT 23.485 191.340 23.845 191.920 ;
        RECT 24.025 191.590 24.275 192.090 ;
        RECT 24.445 191.420 24.785 192.450 ;
        RECT 25.075 192.300 25.245 193.060 ;
        RECT 25.460 192.470 25.790 193.230 ;
        RECT 25.075 192.130 25.790 192.300 ;
        RECT 25.960 192.155 26.215 193.060 ;
        RECT 24.985 191.580 25.340 191.950 ;
        RECT 25.620 191.920 25.790 192.130 ;
        RECT 25.620 191.590 25.875 191.920 ;
        RECT 24.100 191.250 24.785 191.420 ;
        RECT 25.620 191.400 25.790 191.590 ;
        RECT 26.045 191.425 26.215 192.155 ;
        RECT 26.390 192.080 26.650 193.230 ;
        RECT 26.825 192.065 27.115 193.230 ;
        RECT 27.285 192.380 27.545 193.060 ;
        RECT 27.715 192.450 27.965 193.230 ;
        RECT 28.215 192.680 28.465 193.060 ;
        RECT 28.635 192.850 28.990 193.230 ;
        RECT 29.995 192.840 30.330 193.060 ;
        RECT 29.595 192.680 29.825 192.720 ;
        RECT 28.215 192.480 29.825 192.680 ;
        RECT 28.215 192.470 29.050 192.480 ;
        RECT 29.640 192.390 29.825 192.480 ;
        RECT 23.145 190.850 23.405 191.180 ;
        RECT 23.615 190.680 23.890 191.160 ;
        RECT 24.100 190.850 24.305 191.250 ;
        RECT 25.075 191.230 25.790 191.400 ;
        RECT 24.475 190.680 24.810 191.080 ;
        RECT 25.075 190.850 25.245 191.230 ;
        RECT 25.460 190.680 25.790 191.060 ;
        RECT 25.960 190.850 26.215 191.425 ;
        RECT 26.390 190.680 26.650 191.520 ;
        RECT 26.825 190.680 27.115 191.405 ;
        RECT 27.285 191.180 27.455 192.380 ;
        RECT 29.155 192.280 29.485 192.310 ;
        RECT 27.685 192.220 29.485 192.280 ;
        RECT 30.075 192.220 30.330 192.840 ;
        RECT 27.625 192.110 30.330 192.220 ;
        RECT 27.625 192.075 27.825 192.110 ;
        RECT 27.625 191.500 27.795 192.075 ;
        RECT 29.155 192.050 30.330 192.110 ;
        RECT 30.510 192.080 30.770 193.230 ;
        RECT 30.945 192.155 31.200 193.060 ;
        RECT 31.370 192.470 31.700 193.230 ;
        RECT 31.915 192.300 32.085 193.060 ;
        RECT 28.025 191.635 28.435 191.940 ;
        RECT 28.605 191.670 28.935 191.880 ;
        RECT 27.625 191.380 27.895 191.500 ;
        RECT 27.625 191.335 28.470 191.380 ;
        RECT 27.715 191.210 28.470 191.335 ;
        RECT 28.725 191.270 28.935 191.670 ;
        RECT 29.180 191.670 29.655 191.880 ;
        RECT 29.845 191.670 30.335 191.870 ;
        RECT 29.180 191.270 29.400 191.670 ;
        RECT 27.285 190.850 27.545 191.180 ;
        RECT 28.300 191.060 28.470 191.210 ;
        RECT 27.715 190.680 28.045 191.040 ;
        RECT 28.300 190.850 29.600 191.060 ;
        RECT 29.875 190.680 30.330 191.445 ;
        RECT 30.510 190.680 30.770 191.520 ;
        RECT 30.945 191.425 31.115 192.155 ;
        RECT 31.370 192.130 32.085 192.300 ;
        RECT 31.370 191.920 31.540 192.130 ;
        RECT 32.350 192.080 32.610 193.230 ;
        RECT 32.785 192.155 33.040 193.060 ;
        RECT 33.210 192.470 33.540 193.230 ;
        RECT 33.755 192.300 33.925 193.060 ;
        RECT 31.285 191.590 31.540 191.920 ;
        RECT 30.945 190.850 31.200 191.425 ;
        RECT 31.370 191.400 31.540 191.590 ;
        RECT 31.820 191.580 32.175 191.950 ;
        RECT 31.370 191.230 32.085 191.400 ;
        RECT 31.370 190.680 31.700 191.060 ;
        RECT 31.915 190.850 32.085 191.230 ;
        RECT 32.350 190.680 32.610 191.520 ;
        RECT 32.785 191.425 32.955 192.155 ;
        RECT 33.210 192.130 33.925 192.300 ;
        RECT 33.210 191.920 33.380 192.130 ;
        RECT 34.185 192.090 34.445 193.230 ;
        RECT 34.685 192.720 36.300 193.050 ;
        RECT 33.125 191.590 33.380 191.920 ;
        RECT 32.785 190.850 33.040 191.425 ;
        RECT 33.210 191.400 33.380 191.590 ;
        RECT 33.660 191.580 34.015 191.950 ;
        RECT 34.695 191.920 34.865 192.480 ;
        RECT 35.125 192.380 36.300 192.550 ;
        RECT 36.470 192.430 36.750 193.230 ;
        RECT 35.125 192.090 35.455 192.380 ;
        RECT 36.130 192.260 36.300 192.380 ;
        RECT 35.625 191.920 35.870 192.210 ;
        RECT 36.130 192.090 36.790 192.260 ;
        RECT 36.960 192.090 37.235 193.060 ;
        RECT 36.620 191.920 36.790 192.090 ;
        RECT 34.190 191.670 34.525 191.920 ;
        RECT 34.695 191.590 35.410 191.920 ;
        RECT 35.625 191.590 36.450 191.920 ;
        RECT 36.620 191.590 36.895 191.920 ;
        RECT 34.695 191.500 34.945 191.590 ;
        RECT 33.210 191.230 33.925 191.400 ;
        RECT 33.210 190.680 33.540 191.060 ;
        RECT 33.755 190.850 33.925 191.230 ;
        RECT 34.185 190.680 34.445 191.500 ;
        RECT 34.615 191.080 34.945 191.500 ;
        RECT 36.620 191.420 36.790 191.590 ;
        RECT 35.125 191.250 36.790 191.420 ;
        RECT 37.065 191.355 37.235 192.090 ;
        RECT 37.410 192.080 37.670 193.230 ;
        RECT 37.845 192.155 38.100 193.060 ;
        RECT 38.270 192.470 38.600 193.230 ;
        RECT 38.815 192.300 38.985 193.060 ;
        RECT 35.125 190.850 35.385 191.250 ;
        RECT 35.555 190.680 35.885 191.080 ;
        RECT 36.055 190.900 36.225 191.250 ;
        RECT 36.395 190.680 36.770 191.080 ;
        RECT 36.960 191.010 37.235 191.355 ;
        RECT 37.410 190.680 37.670 191.520 ;
        RECT 37.845 191.425 38.015 192.155 ;
        RECT 38.270 192.130 38.985 192.300 ;
        RECT 38.270 191.920 38.440 192.130 ;
        RECT 39.705 192.065 39.995 193.230 ;
        RECT 40.165 192.155 40.435 193.060 ;
        RECT 40.605 192.470 40.935 193.230 ;
        RECT 41.115 192.300 41.285 193.060 ;
        RECT 38.185 191.590 38.440 191.920 ;
        RECT 37.845 190.850 38.100 191.425 ;
        RECT 38.270 191.400 38.440 191.590 ;
        RECT 38.720 191.580 39.075 191.950 ;
        RECT 38.270 191.230 38.985 191.400 ;
        RECT 38.270 190.680 38.600 191.060 ;
        RECT 38.815 190.850 38.985 191.230 ;
        RECT 39.705 190.680 39.995 191.405 ;
        RECT 40.165 191.355 40.335 192.155 ;
        RECT 40.620 192.130 41.285 192.300 ;
        RECT 41.635 192.300 41.805 193.060 ;
        RECT 41.985 192.470 42.315 193.230 ;
        RECT 41.635 192.130 42.300 192.300 ;
        RECT 42.485 192.155 42.755 193.060 ;
        RECT 40.620 191.985 40.790 192.130 ;
        RECT 40.505 191.655 40.790 191.985 ;
        RECT 42.130 191.985 42.300 192.130 ;
        RECT 40.620 191.400 40.790 191.655 ;
        RECT 41.025 191.580 41.355 191.950 ;
        RECT 41.565 191.580 41.895 191.950 ;
        RECT 42.130 191.655 42.415 191.985 ;
        RECT 42.130 191.400 42.300 191.655 ;
        RECT 40.165 190.850 40.425 191.355 ;
        RECT 40.620 191.230 41.285 191.400 ;
        RECT 40.605 190.680 40.935 191.060 ;
        RECT 41.115 190.850 41.285 191.230 ;
        RECT 41.635 191.230 42.300 191.400 ;
        RECT 42.585 191.355 42.755 192.155 ;
        RECT 42.935 192.090 43.265 193.230 ;
        RECT 43.795 192.260 44.125 193.045 ;
        RECT 43.445 192.090 44.125 192.260 ;
        RECT 44.395 192.300 44.565 193.060 ;
        RECT 44.780 192.470 45.110 193.230 ;
        RECT 44.395 192.130 45.110 192.300 ;
        RECT 45.280 192.155 45.535 193.060 ;
        RECT 42.925 191.670 43.275 191.920 ;
        RECT 43.445 191.490 43.615 192.090 ;
        RECT 43.785 191.670 44.135 191.920 ;
        RECT 44.305 191.580 44.660 191.950 ;
        RECT 44.940 191.920 45.110 192.130 ;
        RECT 44.940 191.590 45.195 191.920 ;
        RECT 41.635 190.850 41.805 191.230 ;
        RECT 41.985 190.680 42.315 191.060 ;
        RECT 42.495 190.850 42.755 191.355 ;
        RECT 42.935 190.680 43.205 191.490 ;
        RECT 43.375 190.850 43.705 191.490 ;
        RECT 43.875 190.680 44.115 191.490 ;
        RECT 44.940 191.400 45.110 191.590 ;
        RECT 45.365 191.425 45.535 192.155 ;
        RECT 45.710 192.080 45.970 193.230 ;
        RECT 46.875 192.720 47.205 193.230 ;
        RECT 46.145 192.380 48.105 192.550 ;
        RECT 44.395 191.230 45.110 191.400 ;
        RECT 44.395 190.850 44.565 191.230 ;
        RECT 44.780 190.680 45.110 191.060 ;
        RECT 45.280 190.850 45.535 191.425 ;
        RECT 45.710 190.680 45.970 191.520 ;
        RECT 46.145 191.420 46.315 192.380 ;
        RECT 46.485 191.590 46.835 192.210 ;
        RECT 47.005 191.590 47.345 192.210 ;
        RECT 47.515 191.590 47.755 192.210 ;
        RECT 47.935 191.840 48.105 192.380 ;
        RECT 48.275 192.040 48.735 193.050 ;
        RECT 48.910 192.840 49.245 193.060 ;
        RECT 50.250 192.850 50.605 193.230 ;
        RECT 48.910 192.220 49.165 192.840 ;
        RECT 49.415 192.680 49.645 192.720 ;
        RECT 50.775 192.680 51.025 193.060 ;
        RECT 49.415 192.480 51.025 192.680 ;
        RECT 49.415 192.390 49.600 192.480 ;
        RECT 50.190 192.470 51.025 192.480 ;
        RECT 51.275 192.450 51.525 193.230 ;
        RECT 51.695 192.380 51.955 193.060 ;
        RECT 49.755 192.280 50.085 192.310 ;
        RECT 49.755 192.220 51.555 192.280 ;
        RECT 48.910 192.110 51.615 192.220 ;
        RECT 48.910 192.050 50.085 192.110 ;
        RECT 51.415 192.075 51.615 192.110 ;
        RECT 47.935 191.670 48.395 191.840 ;
        RECT 48.565 191.420 48.735 192.040 ;
        RECT 48.905 191.670 49.395 191.870 ;
        RECT 49.585 191.670 50.060 191.880 ;
        RECT 46.145 191.250 46.640 191.420 ;
        RECT 46.470 191.000 46.640 191.250 ;
        RECT 46.875 190.680 47.205 191.420 ;
        RECT 47.375 191.250 48.735 191.420 ;
        RECT 47.375 190.905 47.545 191.250 ;
        RECT 47.715 190.680 48.045 191.080 ;
        RECT 48.215 190.850 48.735 191.250 ;
        RECT 48.910 190.680 49.365 191.445 ;
        RECT 49.840 191.270 50.060 191.670 ;
        RECT 50.305 191.670 50.635 191.880 ;
        RECT 50.305 191.270 50.515 191.670 ;
        RECT 50.805 191.635 51.215 191.940 ;
        RECT 51.445 191.500 51.615 192.075 ;
        RECT 51.345 191.380 51.615 191.500 ;
        RECT 50.770 191.335 51.615 191.380 ;
        RECT 50.770 191.210 51.525 191.335 ;
        RECT 50.770 191.060 50.940 191.210 ;
        RECT 51.785 191.190 51.955 192.380 ;
        RECT 52.585 192.065 52.875 193.230 ;
        RECT 53.975 192.090 54.305 193.230 ;
        RECT 54.835 192.260 55.165 193.045 ;
        RECT 54.485 192.090 55.165 192.260 ;
        RECT 53.965 191.670 54.315 191.920 ;
        RECT 54.485 191.490 54.655 192.090 ;
        RECT 55.805 192.040 56.265 193.050 ;
        RECT 57.335 192.720 57.665 193.230 ;
        RECT 56.435 192.380 58.395 192.550 ;
        RECT 54.825 191.670 55.175 191.920 ;
        RECT 51.725 191.180 51.955 191.190 ;
        RECT 49.640 190.850 50.940 191.060 ;
        RECT 51.195 190.680 51.525 191.040 ;
        RECT 51.695 190.850 51.955 191.180 ;
        RECT 52.585 190.680 52.875 191.405 ;
        RECT 53.975 190.680 54.245 191.490 ;
        RECT 54.415 190.850 54.745 191.490 ;
        RECT 54.915 190.680 55.155 191.490 ;
        RECT 55.805 191.420 55.975 192.040 ;
        RECT 56.435 191.840 56.605 192.380 ;
        RECT 56.145 191.670 56.605 191.840 ;
        RECT 56.785 191.590 57.025 192.210 ;
        RECT 57.195 191.590 57.535 192.210 ;
        RECT 57.705 191.590 58.055 192.210 ;
        RECT 58.225 191.420 58.395 192.380 ;
        RECT 58.655 192.300 58.825 193.060 ;
        RECT 59.040 192.470 59.370 193.230 ;
        RECT 58.655 192.130 59.370 192.300 ;
        RECT 59.540 192.155 59.795 193.060 ;
        RECT 58.565 191.580 58.920 191.950 ;
        RECT 59.200 191.920 59.370 192.130 ;
        RECT 59.200 191.590 59.455 191.920 ;
        RECT 55.805 191.250 57.165 191.420 ;
        RECT 55.805 190.850 56.325 191.250 ;
        RECT 56.495 190.680 56.825 191.080 ;
        RECT 56.995 190.905 57.165 191.250 ;
        RECT 57.335 190.680 57.665 191.420 ;
        RECT 57.900 191.250 58.395 191.420 ;
        RECT 59.200 191.400 59.370 191.590 ;
        RECT 59.625 191.425 59.795 192.155 ;
        RECT 59.970 192.080 60.230 193.230 ;
        RECT 60.405 192.155 60.675 193.060 ;
        RECT 60.845 192.470 61.175 193.230 ;
        RECT 61.355 192.300 61.525 193.060 ;
        RECT 57.900 191.000 58.070 191.250 ;
        RECT 58.655 191.230 59.370 191.400 ;
        RECT 58.655 190.850 58.825 191.230 ;
        RECT 59.040 190.680 59.370 191.060 ;
        RECT 59.540 190.850 59.795 191.425 ;
        RECT 59.970 190.680 60.230 191.520 ;
        RECT 60.405 191.355 60.575 192.155 ;
        RECT 60.860 192.130 61.525 192.300 ;
        RECT 61.795 192.260 62.125 193.045 ;
        RECT 60.860 191.985 61.030 192.130 ;
        RECT 61.795 192.090 62.475 192.260 ;
        RECT 62.655 192.090 62.985 193.230 ;
        RECT 63.175 192.090 63.505 193.230 ;
        RECT 64.035 192.260 64.365 193.045 ;
        RECT 63.685 192.090 64.365 192.260 ;
        RECT 60.745 191.655 61.030 191.985 ;
        RECT 60.860 191.400 61.030 191.655 ;
        RECT 61.265 191.580 61.595 191.950 ;
        RECT 61.785 191.670 62.135 191.920 ;
        RECT 62.305 191.490 62.475 192.090 ;
        RECT 62.645 191.670 62.995 191.920 ;
        RECT 63.165 191.670 63.515 191.920 ;
        RECT 63.685 191.490 63.855 192.090 ;
        RECT 65.465 192.065 65.755 193.230 ;
        RECT 66.015 192.300 66.185 193.060 ;
        RECT 66.400 192.470 66.730 193.230 ;
        RECT 66.015 192.130 66.730 192.300 ;
        RECT 66.900 192.155 67.155 193.060 ;
        RECT 64.025 191.670 64.375 191.920 ;
        RECT 65.925 191.580 66.280 191.950 ;
        RECT 66.560 191.920 66.730 192.130 ;
        RECT 66.560 191.590 66.815 191.920 ;
        RECT 60.405 190.850 60.665 191.355 ;
        RECT 60.860 191.230 61.525 191.400 ;
        RECT 60.845 190.680 61.175 191.060 ;
        RECT 61.355 190.850 61.525 191.230 ;
        RECT 61.805 190.680 62.045 191.490 ;
        RECT 62.215 190.850 62.545 191.490 ;
        RECT 62.715 190.680 62.985 191.490 ;
        RECT 63.175 190.680 63.445 191.490 ;
        RECT 63.615 190.850 63.945 191.490 ;
        RECT 64.115 190.680 64.355 191.490 ;
        RECT 65.465 190.680 65.755 191.405 ;
        RECT 66.560 191.400 66.730 191.590 ;
        RECT 66.985 191.425 67.155 192.155 ;
        RECT 67.330 192.080 67.590 193.230 ;
        RECT 67.765 192.140 69.435 193.230 ;
        RECT 66.015 191.230 66.730 191.400 ;
        RECT 66.015 190.850 66.185 191.230 ;
        RECT 66.400 190.680 66.730 191.060 ;
        RECT 66.900 190.850 67.155 191.425 ;
        RECT 67.330 190.680 67.590 191.520 ;
        RECT 67.765 191.450 68.515 191.970 ;
        RECT 68.685 191.620 69.435 192.140 ;
        RECT 69.695 192.300 69.865 193.060 ;
        RECT 70.045 192.470 70.375 193.230 ;
        RECT 69.695 192.130 70.360 192.300 ;
        RECT 70.545 192.155 70.815 193.060 ;
        RECT 70.190 191.985 70.360 192.130 ;
        RECT 69.625 191.580 69.955 191.950 ;
        RECT 70.190 191.655 70.475 191.985 ;
        RECT 67.765 190.680 69.435 191.450 ;
        RECT 70.190 191.400 70.360 191.655 ;
        RECT 69.695 191.230 70.360 191.400 ;
        RECT 70.645 191.355 70.815 192.155 ;
        RECT 70.995 192.090 71.325 193.230 ;
        RECT 71.855 192.260 72.185 193.045 ;
        RECT 71.505 192.090 72.185 192.260 ;
        RECT 72.455 192.300 72.625 193.060 ;
        RECT 72.805 192.470 73.135 193.230 ;
        RECT 72.455 192.130 73.120 192.300 ;
        RECT 73.305 192.155 73.575 193.060 ;
        RECT 70.985 191.670 71.335 191.920 ;
        RECT 71.505 191.490 71.675 192.090 ;
        RECT 72.950 191.985 73.120 192.130 ;
        RECT 71.845 191.670 72.195 191.920 ;
        RECT 72.385 191.580 72.715 191.950 ;
        RECT 72.950 191.655 73.235 191.985 ;
        RECT 69.695 190.850 69.865 191.230 ;
        RECT 70.045 190.680 70.375 191.060 ;
        RECT 70.555 190.850 70.815 191.355 ;
        RECT 70.995 190.680 71.265 191.490 ;
        RECT 71.435 190.850 71.765 191.490 ;
        RECT 71.935 190.680 72.175 191.490 ;
        RECT 72.950 191.400 73.120 191.655 ;
        RECT 72.455 191.230 73.120 191.400 ;
        RECT 73.405 191.355 73.575 192.155 ;
        RECT 73.835 192.300 74.005 193.060 ;
        RECT 74.220 192.470 74.550 193.230 ;
        RECT 73.835 192.130 74.550 192.300 ;
        RECT 74.720 192.155 74.975 193.060 ;
        RECT 73.745 191.580 74.100 191.950 ;
        RECT 74.380 191.920 74.550 192.130 ;
        RECT 74.380 191.590 74.635 191.920 ;
        RECT 74.380 191.400 74.550 191.590 ;
        RECT 74.805 191.425 74.975 192.155 ;
        RECT 75.150 192.080 75.410 193.230 ;
        RECT 75.585 192.040 76.045 193.050 ;
        RECT 77.115 192.720 77.445 193.230 ;
        RECT 76.215 192.380 78.175 192.550 ;
        RECT 72.455 190.850 72.625 191.230 ;
        RECT 72.805 190.680 73.135 191.060 ;
        RECT 73.315 190.850 73.575 191.355 ;
        RECT 73.835 191.230 74.550 191.400 ;
        RECT 73.835 190.850 74.005 191.230 ;
        RECT 74.220 190.680 74.550 191.060 ;
        RECT 74.720 190.850 74.975 191.425 ;
        RECT 75.150 190.680 75.410 191.520 ;
        RECT 75.585 191.420 75.755 192.040 ;
        RECT 76.215 191.840 76.385 192.380 ;
        RECT 75.925 191.670 76.385 191.840 ;
        RECT 76.565 191.590 76.805 192.210 ;
        RECT 76.975 191.590 77.315 192.210 ;
        RECT 77.485 191.590 77.835 192.210 ;
        RECT 78.005 191.420 78.175 192.380 ;
        RECT 78.345 192.065 78.635 193.230 ;
        RECT 78.810 192.840 79.145 193.060 ;
        RECT 80.150 192.850 80.505 193.230 ;
        RECT 78.810 192.220 79.065 192.840 ;
        RECT 79.315 192.680 79.545 192.720 ;
        RECT 80.675 192.680 80.925 193.060 ;
        RECT 79.315 192.480 80.925 192.680 ;
        RECT 79.315 192.390 79.500 192.480 ;
        RECT 80.090 192.470 80.925 192.480 ;
        RECT 81.175 192.450 81.425 193.230 ;
        RECT 81.595 192.380 81.855 193.060 ;
        RECT 79.655 192.280 79.985 192.310 ;
        RECT 79.655 192.220 81.455 192.280 ;
        RECT 78.810 192.110 81.515 192.220 ;
        RECT 78.810 192.050 79.985 192.110 ;
        RECT 81.315 192.075 81.515 192.110 ;
        RECT 78.805 191.670 79.295 191.870 ;
        RECT 79.485 191.670 79.960 191.880 ;
        RECT 75.585 191.250 76.945 191.420 ;
        RECT 75.585 190.850 76.105 191.250 ;
        RECT 76.275 190.680 76.605 191.080 ;
        RECT 76.775 190.905 76.945 191.250 ;
        RECT 77.115 190.680 77.445 191.420 ;
        RECT 77.680 191.250 78.175 191.420 ;
        RECT 77.680 191.000 77.850 191.250 ;
        RECT 78.345 190.680 78.635 191.405 ;
        RECT 78.810 190.680 79.265 191.445 ;
        RECT 79.740 191.270 79.960 191.670 ;
        RECT 80.205 191.670 80.535 191.880 ;
        RECT 80.205 191.270 80.415 191.670 ;
        RECT 80.705 191.635 81.115 191.940 ;
        RECT 81.345 191.500 81.515 192.075 ;
        RECT 81.245 191.380 81.515 191.500 ;
        RECT 80.670 191.335 81.515 191.380 ;
        RECT 80.670 191.210 81.425 191.335 ;
        RECT 80.670 191.060 80.840 191.210 ;
        RECT 81.685 191.180 81.855 192.380 ;
        RECT 82.035 192.090 82.365 193.230 ;
        RECT 82.895 192.260 83.225 193.045 ;
        RECT 82.545 192.090 83.225 192.260 ;
        RECT 83.495 192.300 83.665 193.060 ;
        RECT 83.880 192.470 84.210 193.230 ;
        RECT 83.495 192.130 84.210 192.300 ;
        RECT 84.380 192.155 84.635 193.060 ;
        RECT 82.025 191.670 82.375 191.920 ;
        RECT 82.545 191.490 82.715 192.090 ;
        RECT 82.885 191.670 83.235 191.920 ;
        RECT 83.405 191.580 83.760 191.950 ;
        RECT 84.040 191.920 84.210 192.130 ;
        RECT 84.040 191.590 84.295 191.920 ;
        RECT 79.540 190.850 80.840 191.060 ;
        RECT 81.095 190.680 81.425 191.040 ;
        RECT 81.595 190.850 81.855 191.180 ;
        RECT 82.035 190.680 82.305 191.490 ;
        RECT 82.475 190.850 82.805 191.490 ;
        RECT 82.975 190.680 83.215 191.490 ;
        RECT 84.040 191.400 84.210 191.590 ;
        RECT 84.465 191.425 84.635 192.155 ;
        RECT 84.810 192.080 85.070 193.230 ;
        RECT 86.165 192.155 86.435 193.060 ;
        RECT 86.605 192.470 86.935 193.230 ;
        RECT 87.115 192.300 87.285 193.060 ;
        RECT 83.495 191.230 84.210 191.400 ;
        RECT 83.495 190.850 83.665 191.230 ;
        RECT 83.880 190.680 84.210 191.060 ;
        RECT 84.380 190.850 84.635 191.425 ;
        RECT 84.810 190.680 85.070 191.520 ;
        RECT 86.165 191.355 86.335 192.155 ;
        RECT 86.620 192.130 87.285 192.300 ;
        RECT 87.550 192.840 87.885 193.060 ;
        RECT 88.890 192.850 89.245 193.230 ;
        RECT 87.550 192.220 87.805 192.840 ;
        RECT 88.055 192.680 88.285 192.720 ;
        RECT 89.415 192.680 89.665 193.060 ;
        RECT 88.055 192.480 89.665 192.680 ;
        RECT 88.055 192.390 88.240 192.480 ;
        RECT 88.830 192.470 89.665 192.480 ;
        RECT 89.915 192.450 90.165 193.230 ;
        RECT 90.335 192.380 90.595 193.060 ;
        RECT 88.395 192.280 88.725 192.310 ;
        RECT 88.395 192.220 90.195 192.280 ;
        RECT 86.620 191.985 86.790 192.130 ;
        RECT 87.550 192.110 90.255 192.220 ;
        RECT 87.550 192.050 88.725 192.110 ;
        RECT 90.055 192.075 90.255 192.110 ;
        RECT 86.505 191.655 86.790 191.985 ;
        RECT 86.620 191.400 86.790 191.655 ;
        RECT 87.025 191.580 87.355 191.950 ;
        RECT 87.545 191.670 88.035 191.870 ;
        RECT 88.225 191.670 88.700 191.880 ;
        RECT 86.165 190.850 86.425 191.355 ;
        RECT 86.620 191.230 87.285 191.400 ;
        RECT 86.605 190.680 86.935 191.060 ;
        RECT 87.115 190.850 87.285 191.230 ;
        RECT 87.550 190.680 88.005 191.445 ;
        RECT 88.480 191.270 88.700 191.670 ;
        RECT 88.945 191.670 89.275 191.880 ;
        RECT 88.945 191.270 89.155 191.670 ;
        RECT 89.445 191.635 89.855 191.940 ;
        RECT 90.085 191.500 90.255 192.075 ;
        RECT 89.985 191.380 90.255 191.500 ;
        RECT 89.410 191.335 90.255 191.380 ;
        RECT 89.410 191.210 90.165 191.335 ;
        RECT 89.410 191.060 89.580 191.210 ;
        RECT 90.425 191.180 90.595 192.380 ;
        RECT 91.225 192.065 91.515 193.230 ;
        RECT 92.695 192.300 92.865 193.060 ;
        RECT 93.080 192.470 93.410 193.230 ;
        RECT 92.695 192.130 93.410 192.300 ;
        RECT 93.580 192.155 93.835 193.060 ;
        RECT 92.605 191.580 92.960 191.950 ;
        RECT 93.240 191.920 93.410 192.130 ;
        RECT 93.240 191.590 93.495 191.920 ;
        RECT 88.280 190.850 89.580 191.060 ;
        RECT 89.835 190.680 90.165 191.040 ;
        RECT 90.335 190.850 90.595 191.180 ;
        RECT 91.225 190.680 91.515 191.405 ;
        RECT 93.240 191.400 93.410 191.590 ;
        RECT 93.665 191.425 93.835 192.155 ;
        RECT 94.010 192.080 94.270 193.230 ;
        RECT 95.635 192.720 95.965 193.230 ;
        RECT 94.905 192.380 96.865 192.550 ;
        RECT 92.695 191.230 93.410 191.400 ;
        RECT 92.695 190.850 92.865 191.230 ;
        RECT 93.080 190.680 93.410 191.060 ;
        RECT 93.580 190.850 93.835 191.425 ;
        RECT 94.010 190.680 94.270 191.520 ;
        RECT 94.905 191.420 95.075 192.380 ;
        RECT 95.245 191.590 95.595 192.210 ;
        RECT 95.765 191.590 96.105 192.210 ;
        RECT 96.275 191.590 96.515 192.210 ;
        RECT 96.695 191.840 96.865 192.380 ;
        RECT 97.035 192.040 97.495 193.050 ;
        RECT 97.670 192.840 98.005 193.060 ;
        RECT 99.010 192.850 99.365 193.230 ;
        RECT 97.670 192.220 97.925 192.840 ;
        RECT 98.175 192.680 98.405 192.720 ;
        RECT 99.535 192.680 99.785 193.060 ;
        RECT 98.175 192.480 99.785 192.680 ;
        RECT 98.175 192.390 98.360 192.480 ;
        RECT 98.950 192.470 99.785 192.480 ;
        RECT 100.035 192.450 100.285 193.230 ;
        RECT 100.455 192.380 100.715 193.060 ;
        RECT 98.515 192.280 98.845 192.310 ;
        RECT 98.515 192.220 100.315 192.280 ;
        RECT 97.670 192.110 100.375 192.220 ;
        RECT 97.670 192.050 98.845 192.110 ;
        RECT 100.175 192.075 100.375 192.110 ;
        RECT 96.695 191.670 97.155 191.840 ;
        RECT 97.325 191.420 97.495 192.040 ;
        RECT 97.665 191.670 98.155 191.870 ;
        RECT 98.345 191.670 98.820 191.880 ;
        RECT 94.905 191.250 95.400 191.420 ;
        RECT 95.230 191.000 95.400 191.250 ;
        RECT 95.635 190.680 95.965 191.420 ;
        RECT 96.135 191.250 97.495 191.420 ;
        RECT 96.135 190.905 96.305 191.250 ;
        RECT 96.475 190.680 96.805 191.080 ;
        RECT 96.975 190.850 97.495 191.250 ;
        RECT 97.670 190.680 98.125 191.445 ;
        RECT 98.600 191.270 98.820 191.670 ;
        RECT 99.065 191.670 99.395 191.880 ;
        RECT 99.065 191.270 99.275 191.670 ;
        RECT 99.565 191.635 99.975 191.940 ;
        RECT 100.205 191.500 100.375 192.075 ;
        RECT 100.105 191.380 100.375 191.500 ;
        RECT 99.530 191.335 100.375 191.380 ;
        RECT 99.530 191.210 100.285 191.335 ;
        RECT 99.530 191.060 99.700 191.210 ;
        RECT 100.545 191.190 100.715 192.380 ;
        RECT 101.810 192.080 102.070 193.230 ;
        RECT 102.245 192.155 102.500 193.060 ;
        RECT 102.670 192.470 103.000 193.230 ;
        RECT 103.215 192.300 103.385 193.060 ;
        RECT 100.485 191.180 100.715 191.190 ;
        RECT 98.400 190.850 99.700 191.060 ;
        RECT 99.955 190.680 100.285 191.040 ;
        RECT 100.455 190.850 100.715 191.180 ;
        RECT 101.810 190.680 102.070 191.520 ;
        RECT 102.245 191.425 102.415 192.155 ;
        RECT 102.670 192.130 103.385 192.300 ;
        RECT 102.670 191.920 102.840 192.130 ;
        RECT 104.105 192.065 104.395 193.230 ;
        RECT 104.875 192.390 105.045 193.230 ;
        RECT 105.255 192.220 105.505 193.060 ;
        RECT 105.715 192.390 105.885 193.230 ;
        RECT 106.055 192.220 106.345 193.060 ;
        RECT 104.620 192.050 106.345 192.220 ;
        RECT 106.555 192.170 106.725 193.230 ;
        RECT 107.020 192.850 107.350 193.230 ;
        RECT 107.530 192.680 107.700 192.970 ;
        RECT 107.870 192.770 108.120 193.230 ;
        RECT 106.900 192.510 107.700 192.680 ;
        RECT 108.290 192.720 109.160 193.060 ;
        RECT 102.585 191.590 102.840 191.920 ;
        RECT 102.245 190.850 102.500 191.425 ;
        RECT 102.670 191.400 102.840 191.590 ;
        RECT 103.120 191.580 103.475 191.950 ;
        RECT 104.620 191.500 105.030 192.050 ;
        RECT 106.900 191.890 107.070 192.510 ;
        RECT 108.290 192.340 108.460 192.720 ;
        RECT 109.395 192.600 109.565 193.060 ;
        RECT 109.735 192.770 110.105 193.230 ;
        RECT 110.400 192.630 110.570 192.970 ;
        RECT 110.740 192.800 111.070 193.230 ;
        RECT 111.305 192.630 111.475 192.970 ;
        RECT 107.240 192.170 108.460 192.340 ;
        RECT 108.630 192.260 109.090 192.550 ;
        RECT 109.395 192.430 109.955 192.600 ;
        RECT 110.400 192.460 111.475 192.630 ;
        RECT 111.645 192.730 112.325 193.060 ;
        RECT 112.540 192.730 112.790 193.060 ;
        RECT 112.960 192.770 113.210 193.230 ;
        RECT 109.785 192.290 109.955 192.430 ;
        RECT 108.630 192.250 109.595 192.260 ;
        RECT 108.290 192.080 108.460 192.170 ;
        RECT 108.920 192.090 109.595 192.250 ;
        RECT 106.900 191.880 107.245 191.890 ;
        RECT 105.215 191.670 107.245 191.880 ;
        RECT 102.670 191.230 103.385 191.400 ;
        RECT 102.670 190.680 103.000 191.060 ;
        RECT 103.215 190.850 103.385 191.230 ;
        RECT 104.105 190.680 104.395 191.405 ;
        RECT 104.620 191.330 106.385 191.500 ;
        RECT 104.875 190.680 105.045 191.150 ;
        RECT 105.215 190.850 105.545 191.330 ;
        RECT 105.715 190.680 105.885 191.150 ;
        RECT 106.055 190.850 106.385 191.330 ;
        RECT 106.555 190.680 106.725 191.490 ;
        RECT 106.920 191.415 107.245 191.670 ;
        RECT 106.925 191.060 107.245 191.415 ;
        RECT 107.415 191.630 107.955 192.000 ;
        RECT 108.290 191.910 108.695 192.080 ;
        RECT 107.415 191.230 107.655 191.630 ;
        RECT 108.135 191.460 108.355 191.740 ;
        RECT 107.825 191.290 108.355 191.460 ;
        RECT 107.825 191.060 107.995 191.290 ;
        RECT 108.525 191.130 108.695 191.910 ;
        RECT 108.865 191.300 109.215 191.920 ;
        RECT 109.385 191.300 109.595 192.090 ;
        RECT 109.785 192.120 111.285 192.290 ;
        RECT 109.785 191.430 109.955 192.120 ;
        RECT 111.645 191.950 111.815 192.730 ;
        RECT 112.620 192.600 112.790 192.730 ;
        RECT 110.125 191.780 111.815 191.950 ;
        RECT 111.985 192.170 112.450 192.560 ;
        RECT 112.620 192.430 113.015 192.600 ;
        RECT 110.125 191.600 110.295 191.780 ;
        RECT 106.925 190.890 107.995 191.060 ;
        RECT 108.165 190.680 108.355 191.120 ;
        RECT 108.525 190.850 109.475 191.130 ;
        RECT 109.785 191.040 110.045 191.430 ;
        RECT 110.465 191.360 111.255 191.610 ;
        RECT 109.695 190.870 110.045 191.040 ;
        RECT 110.255 190.680 110.585 191.140 ;
        RECT 111.460 191.070 111.630 191.780 ;
        RECT 111.985 191.580 112.155 192.170 ;
        RECT 111.800 191.360 112.155 191.580 ;
        RECT 112.325 191.360 112.675 191.980 ;
        RECT 112.845 191.070 113.015 192.430 ;
        RECT 113.380 192.260 113.705 193.045 ;
        RECT 113.185 191.210 113.645 192.260 ;
        RECT 111.460 190.900 112.315 191.070 ;
        RECT 112.520 190.900 113.015 191.070 ;
        RECT 113.185 190.680 113.515 191.040 ;
        RECT 113.875 190.940 114.045 193.060 ;
        RECT 114.215 192.730 114.545 193.230 ;
        RECT 114.715 192.560 114.970 193.060 ;
        RECT 114.220 192.390 114.970 192.560 ;
        RECT 114.220 191.400 114.450 192.390 ;
        RECT 114.620 191.570 114.970 192.220 ;
        RECT 115.150 192.080 115.410 193.230 ;
        RECT 115.585 192.155 115.840 193.060 ;
        RECT 116.010 192.470 116.340 193.230 ;
        RECT 116.555 192.300 116.725 193.060 ;
        RECT 114.220 191.230 114.970 191.400 ;
        RECT 114.215 190.680 114.545 191.060 ;
        RECT 114.715 190.940 114.970 191.230 ;
        RECT 115.150 190.680 115.410 191.520 ;
        RECT 115.585 191.425 115.755 192.155 ;
        RECT 116.010 192.130 116.725 192.300 ;
        RECT 116.010 191.920 116.180 192.130 ;
        RECT 116.985 192.065 117.275 193.230 ;
        RECT 117.535 192.300 117.705 193.060 ;
        RECT 117.885 192.470 118.215 193.230 ;
        RECT 117.535 192.130 118.200 192.300 ;
        RECT 118.385 192.155 118.655 193.060 ;
        RECT 118.030 191.985 118.200 192.130 ;
        RECT 115.925 191.590 116.180 191.920 ;
        RECT 115.585 190.850 115.840 191.425 ;
        RECT 116.010 191.400 116.180 191.590 ;
        RECT 116.460 191.580 116.815 191.950 ;
        RECT 117.465 191.580 117.795 191.950 ;
        RECT 118.030 191.655 118.315 191.985 ;
        RECT 116.010 191.230 116.725 191.400 ;
        RECT 116.010 190.680 116.340 191.060 ;
        RECT 116.555 190.850 116.725 191.230 ;
        RECT 116.985 190.680 117.275 191.405 ;
        RECT 118.030 191.400 118.200 191.655 ;
        RECT 117.535 191.230 118.200 191.400 ;
        RECT 118.485 191.355 118.655 192.155 ;
        RECT 117.535 190.850 117.705 191.230 ;
        RECT 117.885 190.680 118.215 191.060 ;
        RECT 118.395 190.850 118.655 191.355 ;
        RECT 119.750 192.510 120.085 193.020 ;
        RECT 119.750 191.155 120.005 192.510 ;
        RECT 120.335 192.430 120.665 193.230 ;
        RECT 120.910 192.640 121.195 193.060 ;
        RECT 121.450 192.810 121.780 193.230 ;
        RECT 122.005 192.890 123.165 193.060 ;
        RECT 122.005 192.640 122.335 192.890 ;
        RECT 120.910 192.470 122.335 192.640 ;
        RECT 122.565 192.260 122.735 192.720 ;
        RECT 122.995 192.390 123.165 192.890 ;
        RECT 123.515 192.610 123.685 193.040 ;
        RECT 123.855 192.780 124.185 193.230 ;
        RECT 123.515 192.380 124.190 192.610 ;
        RECT 120.365 192.090 122.735 192.260 ;
        RECT 120.365 191.920 120.535 192.090 ;
        RECT 122.985 191.920 123.190 192.210 ;
        RECT 120.230 191.590 120.535 191.920 ;
        RECT 120.730 191.870 120.980 191.920 ;
        RECT 120.725 191.700 120.980 191.870 ;
        RECT 120.730 191.590 120.980 191.700 ;
        RECT 120.365 191.420 120.535 191.590 ;
        RECT 121.190 191.530 121.460 191.920 ;
        RECT 121.650 191.870 121.940 191.920 ;
        RECT 121.645 191.700 121.940 191.870 ;
        RECT 120.365 191.250 120.925 191.420 ;
        RECT 121.185 191.360 121.460 191.530 ;
        RECT 121.190 191.260 121.460 191.360 ;
        RECT 121.650 191.260 121.940 191.700 ;
        RECT 122.110 191.255 122.530 191.920 ;
        RECT 122.840 191.870 123.190 191.920 ;
        RECT 122.840 191.700 123.195 191.870 ;
        RECT 122.840 191.590 123.190 191.700 ;
        RECT 119.750 190.895 120.085 191.155 ;
        RECT 120.755 191.080 120.925 191.250 ;
        RECT 120.255 190.680 120.585 191.080 ;
        RECT 120.755 190.910 122.370 191.080 ;
        RECT 122.915 190.680 123.245 191.400 ;
        RECT 123.485 191.360 123.785 192.210 ;
        RECT 123.955 191.730 124.190 192.380 ;
        RECT 124.360 192.070 124.645 193.015 ;
        RECT 124.825 192.760 125.510 193.230 ;
        RECT 124.820 192.240 125.515 192.550 ;
        RECT 125.690 192.175 125.995 192.960 ;
        RECT 124.360 191.920 125.220 192.070 ;
        RECT 124.360 191.900 125.645 191.920 ;
        RECT 123.955 191.400 124.490 191.730 ;
        RECT 124.660 191.540 125.645 191.900 ;
        RECT 123.955 191.250 124.175 191.400 ;
        RECT 123.430 190.680 123.765 191.185 ;
        RECT 123.935 190.875 124.175 191.250 ;
        RECT 124.660 191.205 124.830 191.540 ;
        RECT 125.820 191.370 125.995 192.175 ;
        RECT 126.190 192.080 126.450 193.230 ;
        RECT 126.625 192.155 126.880 193.060 ;
        RECT 127.050 192.470 127.380 193.230 ;
        RECT 127.595 192.300 127.765 193.060 ;
        RECT 124.455 191.010 124.830 191.205 ;
        RECT 124.455 190.865 124.625 191.010 ;
        RECT 125.190 190.680 125.585 191.175 ;
        RECT 125.755 190.850 125.995 191.370 ;
        RECT 126.190 190.680 126.450 191.520 ;
        RECT 126.625 191.425 126.795 192.155 ;
        RECT 127.050 192.130 127.765 192.300 ;
        RECT 128.115 192.300 128.285 193.060 ;
        RECT 128.500 192.470 128.830 193.230 ;
        RECT 128.115 192.130 128.830 192.300 ;
        RECT 129.000 192.155 129.255 193.060 ;
        RECT 127.050 191.920 127.220 192.130 ;
        RECT 126.965 191.590 127.220 191.920 ;
        RECT 126.625 190.850 126.880 191.425 ;
        RECT 127.050 191.400 127.220 191.590 ;
        RECT 127.500 191.580 127.855 191.950 ;
        RECT 128.025 191.580 128.380 191.950 ;
        RECT 128.660 191.920 128.830 192.130 ;
        RECT 128.660 191.590 128.915 191.920 ;
        RECT 128.660 191.400 128.830 191.590 ;
        RECT 129.085 191.425 129.255 192.155 ;
        RECT 129.430 192.080 129.690 193.230 ;
        RECT 129.865 192.065 130.155 193.230 ;
        RECT 130.415 192.300 130.585 193.060 ;
        RECT 130.800 192.470 131.130 193.230 ;
        RECT 130.415 192.130 131.130 192.300 ;
        RECT 131.300 192.155 131.555 193.060 ;
        RECT 130.325 191.580 130.680 191.950 ;
        RECT 130.960 191.920 131.130 192.130 ;
        RECT 130.960 191.590 131.215 191.920 ;
        RECT 127.050 191.230 127.765 191.400 ;
        RECT 127.050 190.680 127.380 191.060 ;
        RECT 127.595 190.850 127.765 191.230 ;
        RECT 128.115 191.230 128.830 191.400 ;
        RECT 128.115 190.850 128.285 191.230 ;
        RECT 128.500 190.680 128.830 191.060 ;
        RECT 129.000 190.850 129.255 191.425 ;
        RECT 129.430 190.680 129.690 191.520 ;
        RECT 129.865 190.680 130.155 191.405 ;
        RECT 130.960 191.400 131.130 191.590 ;
        RECT 131.385 191.425 131.555 192.155 ;
        RECT 131.730 192.080 131.990 193.230 ;
        RECT 133.090 192.080 133.350 193.230 ;
        RECT 133.525 192.155 133.780 193.060 ;
        RECT 133.950 192.470 134.280 193.230 ;
        RECT 134.495 192.300 134.665 193.060 ;
        RECT 130.415 191.230 131.130 191.400 ;
        RECT 130.415 190.850 130.585 191.230 ;
        RECT 130.800 190.680 131.130 191.060 ;
        RECT 131.300 190.850 131.555 191.425 ;
        RECT 131.730 190.680 131.990 191.520 ;
        RECT 133.090 190.680 133.350 191.520 ;
        RECT 133.525 191.425 133.695 192.155 ;
        RECT 133.950 192.130 134.665 192.300 ;
        RECT 133.950 191.920 134.120 192.130 ;
        RECT 134.935 192.090 135.265 193.230 ;
        RECT 135.795 192.260 136.125 193.045 ;
        RECT 136.505 192.560 136.785 193.230 ;
        RECT 136.955 192.340 137.255 192.890 ;
        RECT 137.455 192.510 137.785 193.230 ;
        RECT 137.975 192.510 138.435 193.060 ;
        RECT 139.265 192.560 139.545 193.230 ;
        RECT 135.445 192.090 136.125 192.260 ;
        RECT 133.865 191.590 134.120 191.920 ;
        RECT 133.525 190.850 133.780 191.425 ;
        RECT 133.950 191.400 134.120 191.590 ;
        RECT 134.400 191.580 134.755 191.950 ;
        RECT 134.925 191.670 135.275 191.920 ;
        RECT 135.445 191.490 135.615 192.090 ;
        RECT 136.320 191.920 136.585 192.280 ;
        RECT 136.955 192.170 137.895 192.340 ;
        RECT 137.725 191.920 137.895 192.170 ;
        RECT 135.785 191.670 136.135 191.920 ;
        RECT 136.320 191.670 136.995 191.920 ;
        RECT 137.215 191.670 137.555 191.920 ;
        RECT 137.725 191.590 138.015 191.920 ;
        RECT 137.725 191.500 137.895 191.590 ;
        RECT 133.950 191.230 134.665 191.400 ;
        RECT 133.950 190.680 134.280 191.060 ;
        RECT 134.495 190.850 134.665 191.230 ;
        RECT 134.935 190.680 135.205 191.490 ;
        RECT 135.375 190.850 135.705 191.490 ;
        RECT 135.875 190.680 136.115 191.490 ;
        RECT 136.505 191.310 137.895 191.500 ;
        RECT 136.505 190.950 136.835 191.310 ;
        RECT 138.185 191.140 138.435 192.510 ;
        RECT 139.715 192.340 140.015 192.890 ;
        RECT 140.215 192.510 140.545 193.230 ;
        RECT 140.735 192.510 141.195 193.060 ;
        RECT 139.080 191.920 139.345 192.280 ;
        RECT 139.715 192.170 140.655 192.340 ;
        RECT 140.485 191.920 140.655 192.170 ;
        RECT 139.080 191.670 139.755 191.920 ;
        RECT 139.975 191.670 140.315 191.920 ;
        RECT 140.485 191.590 140.775 191.920 ;
        RECT 140.485 191.500 140.655 191.590 ;
        RECT 137.455 190.680 137.705 191.140 ;
        RECT 137.875 190.850 138.435 191.140 ;
        RECT 139.265 191.310 140.655 191.500 ;
        RECT 139.265 190.950 139.595 191.310 ;
        RECT 140.945 191.140 141.195 192.510 ;
        RECT 141.375 192.260 141.705 193.045 ;
        RECT 141.375 192.090 142.055 192.260 ;
        RECT 142.235 192.090 142.565 193.230 ;
        RECT 141.365 191.670 141.715 191.920 ;
        RECT 141.885 191.490 142.055 192.090 ;
        RECT 142.745 192.065 143.035 193.230 ;
        RECT 143.665 192.260 143.975 193.060 ;
        RECT 144.145 192.430 144.455 193.230 ;
        RECT 144.625 192.600 144.885 193.060 ;
        RECT 145.055 192.770 145.310 193.230 ;
        RECT 145.485 192.600 145.745 193.060 ;
        RECT 144.625 192.430 145.745 192.600 ;
        RECT 143.665 192.090 144.695 192.260 ;
        RECT 142.225 191.670 142.575 191.920 ;
        RECT 140.215 190.680 140.465 191.140 ;
        RECT 140.635 190.850 141.195 191.140 ;
        RECT 141.385 190.680 141.625 191.490 ;
        RECT 141.795 190.850 142.125 191.490 ;
        RECT 142.295 190.680 142.565 191.490 ;
        RECT 142.745 190.680 143.035 191.405 ;
        RECT 143.665 191.180 143.835 192.090 ;
        RECT 144.005 191.350 144.355 191.920 ;
        RECT 144.525 191.840 144.695 192.090 ;
        RECT 145.485 192.180 145.745 192.430 ;
        RECT 145.915 192.360 146.200 193.230 ;
        RECT 145.485 192.010 146.240 192.180 ;
        RECT 144.525 191.670 145.665 191.840 ;
        RECT 145.835 191.500 146.240 192.010 ;
        RECT 146.425 192.140 147.635 193.230 ;
        RECT 146.425 191.600 146.945 192.140 ;
        RECT 144.590 191.330 146.240 191.500 ;
        RECT 147.115 191.430 147.635 191.970 ;
        RECT 143.665 190.850 143.965 191.180 ;
        RECT 144.135 190.680 144.410 191.160 ;
        RECT 144.590 190.940 144.885 191.330 ;
        RECT 145.055 190.680 145.310 191.160 ;
        RECT 145.485 190.940 145.745 191.330 ;
        RECT 145.915 190.680 146.195 191.160 ;
        RECT 146.425 190.680 147.635 191.430 ;
        RECT 13.860 190.510 147.720 190.680 ;
        RECT 109.245 185.185 141.595 185.515 ;
        RECT 109.245 185.015 141.605 185.185 ;
        RECT 8.035 182.490 21.375 182.660 ;
        RECT 8.130 181.960 8.460 182.320 ;
        RECT 8.990 182.130 9.320 182.490 ;
        RECT 9.925 182.130 10.255 182.490 ;
        RECT 9.565 181.960 9.755 182.060 ;
        RECT 10.425 181.960 10.615 182.320 ;
        RECT 10.785 182.130 11.115 182.490 ;
        RECT 8.130 181.770 9.395 181.960 ;
        RECT 8.215 181.580 8.465 181.595 ;
        RECT 8.160 180.960 8.470 181.580 ;
        RECT 8.640 181.250 9.015 181.580 ;
        RECT 9.185 181.555 9.395 181.770 ;
        RECT 9.565 181.730 11.170 181.960 ;
        RECT 9.185 181.220 10.720 181.555 ;
        RECT 9.185 180.995 9.395 181.220 ;
        RECT 10.890 181.040 11.170 181.730 ;
        RECT 11.340 181.720 16.685 182.490 ;
        RECT 16.860 181.740 18.070 182.490 ;
        RECT 18.260 181.980 18.500 182.490 ;
        RECT 11.340 181.200 13.920 181.720 ;
        RECT 8.640 180.825 9.395 180.995 ;
        RECT 8.130 179.940 8.460 180.695 ;
        RECT 8.640 180.110 8.820 180.825 ;
        RECT 9.565 180.815 11.170 181.040 ;
        RECT 14.090 181.030 16.685 181.550 ;
        RECT 16.860 181.200 17.380 181.740 ;
        RECT 17.550 181.030 18.070 181.570 ;
        RECT 18.245 181.250 18.500 181.810 ;
        RECT 18.670 181.750 19.000 182.285 ;
        RECT 19.215 181.750 19.385 182.490 ;
        RECT 19.595 181.840 19.925 182.310 ;
        RECT 20.095 182.010 20.265 182.490 ;
        RECT 20.435 181.840 20.765 182.310 ;
        RECT 20.935 182.010 21.105 182.490 ;
        RECT 18.670 181.080 18.850 181.750 ;
        RECT 19.595 181.670 21.290 181.840 ;
        RECT 19.020 181.250 19.395 181.580 ;
        RECT 19.565 181.330 20.775 181.500 ;
        RECT 19.565 181.080 19.770 181.330 ;
        RECT 20.945 181.080 21.290 181.670 ;
        RECT 9.025 179.940 9.355 180.640 ;
        RECT 9.565 180.110 9.755 180.815 ;
        RECT 10.425 180.810 11.170 180.815 ;
        RECT 9.925 179.940 10.255 180.640 ;
        RECT 10.425 180.110 10.615 180.810 ;
        RECT 10.785 179.940 11.115 180.640 ;
        RECT 11.340 179.940 16.685 181.030 ;
        RECT 16.860 179.940 18.070 181.030 ;
        RECT 18.310 180.910 19.770 181.080 ;
        RECT 20.435 180.910 21.290 181.080 ;
        RECT 47.420 180.940 71.320 181.630 ;
        RECT 71.870 180.940 102.970 181.630 ;
        RECT 18.310 180.110 18.670 180.910 ;
        RECT 20.435 180.740 20.765 180.910 ;
        RECT 47.420 180.770 71.420 180.940 ;
        RECT 19.215 179.940 19.385 180.740 ;
        RECT 19.595 180.570 20.765 180.740 ;
        RECT 19.595 180.110 19.925 180.570 ;
        RECT 20.095 179.940 20.265 180.400 ;
        RECT 20.435 180.110 20.765 180.570 ;
        RECT 20.935 179.940 21.105 180.740 ;
        RECT 8.035 179.770 21.375 179.940 ;
        RECT 34.640 179.840 46.040 180.640 ;
        RECT 8.130 179.015 8.460 179.770 ;
        RECT 8.640 178.885 8.820 179.600 ;
        RECT 9.025 179.070 9.355 179.770 ;
        RECT 9.565 178.895 9.755 179.600 ;
        RECT 9.925 179.070 10.255 179.770 ;
        RECT 10.425 178.900 10.615 179.600 ;
        RECT 10.785 179.070 11.115 179.770 ;
        RECT 11.350 179.015 11.680 179.770 ;
        RECT 10.425 178.895 11.170 178.900 ;
        RECT 8.160 178.130 8.470 178.750 ;
        RECT 8.640 178.715 9.395 178.885 ;
        RECT 9.185 178.490 9.395 178.715 ;
        RECT 9.565 178.670 11.170 178.895 ;
        RECT 11.860 178.885 12.040 179.600 ;
        RECT 12.245 179.070 12.575 179.770 ;
        RECT 12.785 178.895 12.975 179.600 ;
        RECT 13.145 179.070 13.475 179.770 ;
        RECT 13.645 178.900 13.835 179.600 ;
        RECT 14.005 179.070 14.335 179.770 ;
        RECT 13.645 178.895 14.390 178.900 ;
        RECT 8.640 178.130 9.015 178.460 ;
        RECT 9.185 178.155 10.720 178.490 ;
        RECT 9.185 177.940 9.395 178.155 ;
        RECT 10.890 177.980 11.170 178.670 ;
        RECT 11.380 178.130 11.690 178.750 ;
        RECT 11.860 178.715 12.615 178.885 ;
        RECT 12.405 178.490 12.615 178.715 ;
        RECT 12.785 178.670 14.390 178.895 ;
        RECT 11.860 178.130 12.235 178.460 ;
        RECT 12.405 178.155 13.940 178.490 ;
        RECT 8.130 177.750 9.395 177.940 ;
        RECT 9.565 177.750 11.170 177.980 ;
        RECT 12.405 177.940 12.615 178.155 ;
        RECT 14.110 177.980 14.390 178.670 ;
        RECT 14.560 178.605 14.850 179.770 ;
        RECT 15.090 178.800 15.450 179.600 ;
        RECT 15.995 178.970 16.165 179.770 ;
        RECT 16.375 179.140 16.705 179.600 ;
        RECT 16.875 179.310 17.045 179.770 ;
        RECT 17.215 179.140 17.545 179.600 ;
        RECT 16.375 178.970 17.545 179.140 ;
        RECT 17.715 178.970 17.885 179.770 ;
        RECT 17.215 178.800 17.545 178.970 ;
        RECT 18.310 178.800 18.670 179.600 ;
        RECT 19.215 178.970 19.385 179.770 ;
        RECT 19.595 179.140 19.925 179.600 ;
        RECT 20.095 179.310 20.265 179.770 ;
        RECT 20.435 179.140 20.765 179.600 ;
        RECT 19.595 178.970 20.765 179.140 ;
        RECT 20.935 178.970 21.105 179.770 ;
        RECT 35.590 179.755 39.270 179.840 ;
        RECT 35.775 179.295 35.985 179.755 ;
        RECT 20.435 178.800 20.765 178.970 ;
        RECT 36.155 178.805 36.485 179.585 ;
        RECT 36.655 178.955 36.825 179.755 ;
        RECT 15.090 178.630 16.550 178.800 ;
        RECT 17.215 178.630 18.070 178.800 ;
        RECT 18.310 178.630 19.770 178.800 ;
        RECT 20.435 178.630 21.290 178.800 ;
        RECT 15.025 178.415 15.280 178.460 ;
        RECT 15.015 178.165 15.280 178.415 ;
        RECT 11.350 177.750 12.615 177.940 ;
        RECT 12.785 177.750 14.390 177.980 ;
        RECT 8.130 177.390 8.460 177.750 ;
        RECT 9.565 177.650 9.755 177.750 ;
        RECT 8.990 177.220 9.320 177.580 ;
        RECT 9.925 177.220 10.255 177.580 ;
        RECT 10.425 177.390 10.615 177.750 ;
        RECT 10.785 177.220 11.115 177.580 ;
        RECT 11.350 177.390 11.680 177.750 ;
        RECT 12.785 177.650 12.975 177.750 ;
        RECT 12.210 177.220 12.540 177.580 ;
        RECT 13.145 177.220 13.475 177.580 ;
        RECT 13.645 177.390 13.835 177.750 ;
        RECT 14.005 177.220 14.335 177.580 ;
        RECT 14.560 177.220 14.850 177.945 ;
        RECT 15.025 177.900 15.280 178.165 ;
        RECT 15.450 177.960 15.630 178.630 ;
        RECT 15.800 178.130 16.175 178.460 ;
        RECT 16.345 178.380 16.550 178.630 ;
        RECT 16.345 178.210 17.555 178.380 ;
        RECT 17.725 178.040 18.070 178.630 ;
        RECT 15.040 177.220 15.280 177.730 ;
        RECT 15.450 177.425 15.780 177.960 ;
        RECT 15.995 177.220 16.165 177.960 ;
        RECT 16.375 177.870 18.070 178.040 ;
        RECT 18.245 177.900 18.500 178.460 ;
        RECT 18.670 177.960 18.850 178.630 ;
        RECT 19.020 178.130 19.395 178.460 ;
        RECT 19.565 178.380 19.770 178.630 ;
        RECT 19.565 178.210 20.775 178.380 ;
        RECT 20.945 178.040 21.290 178.630 ;
        RECT 35.720 178.785 36.485 178.805 ;
        RECT 36.995 178.785 37.325 179.585 ;
        RECT 35.720 178.615 37.325 178.785 ;
        RECT 37.495 178.615 37.760 179.755 ;
        RECT 35.720 178.440 35.985 178.615 ;
        RECT 38.220 178.605 38.550 179.585 ;
        RECT 38.720 178.615 38.930 179.755 ;
        RECT 39.450 179.720 45.940 179.840 ;
        RECT 35.640 178.140 35.985 178.440 ;
        RECT 36.155 178.440 37.785 178.445 ;
        RECT 38.220 178.440 38.450 178.605 ;
        RECT 36.155 178.195 38.450 178.440 ;
        RECT 38.620 178.195 38.950 178.435 ;
        RECT 37.740 178.190 38.450 178.195 ;
        RECT 16.375 177.400 16.705 177.870 ;
        RECT 16.875 177.220 17.045 177.700 ;
        RECT 17.215 177.400 17.545 177.870 ;
        RECT 17.715 177.220 17.885 177.700 ;
        RECT 18.260 177.220 18.500 177.730 ;
        RECT 18.670 177.425 19.000 177.960 ;
        RECT 19.215 177.220 19.385 177.960 ;
        RECT 19.595 177.870 21.290 178.040 ;
        RECT 35.720 178.025 35.985 178.140 ;
        RECT 19.595 177.400 19.925 177.870 ;
        RECT 20.095 177.220 20.265 177.700 ;
        RECT 20.435 177.400 20.765 177.870 ;
        RECT 35.720 177.845 37.325 178.025 ;
        RECT 20.935 177.220 21.105 177.700 ;
        RECT 8.035 177.050 21.375 177.220 ;
        RECT 35.735 177.205 35.985 177.670 ;
        RECT 36.155 177.375 36.485 177.845 ;
        RECT 36.655 177.205 36.825 177.665 ;
        RECT 36.995 177.375 37.325 177.845 ;
        RECT 38.220 178.005 38.450 178.190 ;
        RECT 37.495 177.205 37.760 177.665 ;
        RECT 38.220 177.375 38.550 178.005 ;
        RECT 38.720 177.205 38.950 178.025 ;
        RECT 39.450 177.240 39.620 179.720 ;
        RECT 40.160 179.210 40.490 179.380 ;
        RECT 40.020 177.955 40.190 178.995 ;
        RECT 40.460 177.955 40.630 178.995 ;
        RECT 40.160 177.570 40.490 177.740 ;
        RECT 41.030 177.240 41.200 179.720 ;
        RECT 41.740 179.210 42.070 179.380 ;
        RECT 8.130 176.520 8.460 176.880 ;
        RECT 8.990 176.690 9.320 177.050 ;
        RECT 9.925 176.690 10.255 177.050 ;
        RECT 9.565 176.520 9.755 176.620 ;
        RECT 10.425 176.520 10.615 176.880 ;
        RECT 10.785 176.690 11.115 177.050 ;
        RECT 11.350 176.520 11.680 176.880 ;
        RECT 12.210 176.690 12.540 177.050 ;
        RECT 13.145 176.690 13.475 177.050 ;
        RECT 12.785 176.520 12.975 176.620 ;
        RECT 13.645 176.520 13.835 176.880 ;
        RECT 14.005 176.690 14.335 177.050 ;
        RECT 8.130 176.330 9.395 176.520 ;
        RECT 8.215 176.140 8.465 176.155 ;
        RECT 8.160 175.520 8.470 176.140 ;
        RECT 8.640 175.810 9.015 176.140 ;
        RECT 9.185 176.115 9.395 176.330 ;
        RECT 9.565 176.290 11.170 176.520 ;
        RECT 11.350 176.330 12.615 176.520 ;
        RECT 9.185 175.780 10.720 176.115 ;
        RECT 9.185 175.555 9.395 175.780 ;
        RECT 10.890 175.600 11.170 176.290 ;
        RECT 8.640 175.385 9.395 175.555 ;
        RECT 8.130 174.500 8.460 175.255 ;
        RECT 8.640 174.670 8.820 175.385 ;
        RECT 9.565 175.375 11.170 175.600 ;
        RECT 11.380 175.520 11.690 176.140 ;
        RECT 11.860 175.810 12.235 176.140 ;
        RECT 12.405 176.115 12.615 176.330 ;
        RECT 12.785 176.290 14.390 176.520 ;
        RECT 14.560 176.325 14.850 177.050 ;
        RECT 15.040 176.540 15.280 177.050 ;
        RECT 12.405 175.780 13.940 176.115 ;
        RECT 12.405 175.555 12.615 175.780 ;
        RECT 14.110 175.600 14.390 176.290 ;
        RECT 15.025 176.105 15.280 176.370 ;
        RECT 15.015 175.855 15.280 176.105 ;
        RECT 15.025 175.810 15.280 175.855 ;
        RECT 15.450 176.310 15.780 176.845 ;
        RECT 15.995 176.310 16.165 177.050 ;
        RECT 16.375 176.400 16.705 176.870 ;
        RECT 16.875 176.570 17.045 177.050 ;
        RECT 17.215 176.400 17.545 176.870 ;
        RECT 17.715 176.570 17.885 177.050 ;
        RECT 18.260 176.540 18.500 177.050 ;
        RECT 9.025 174.500 9.355 175.200 ;
        RECT 9.565 174.670 9.755 175.375 ;
        RECT 10.425 175.370 11.170 175.375 ;
        RECT 11.860 175.385 12.615 175.555 ;
        RECT 9.925 174.500 10.255 175.200 ;
        RECT 10.425 174.670 10.615 175.370 ;
        RECT 10.785 174.500 11.115 175.200 ;
        RECT 11.350 174.500 11.680 175.255 ;
        RECT 11.860 174.670 12.040 175.385 ;
        RECT 12.785 175.375 14.390 175.600 ;
        RECT 12.245 174.500 12.575 175.200 ;
        RECT 12.785 174.670 12.975 175.375 ;
        RECT 13.645 175.370 14.390 175.375 ;
        RECT 13.145 174.500 13.475 175.200 ;
        RECT 13.645 174.670 13.835 175.370 ;
        RECT 14.005 174.500 14.335 175.200 ;
        RECT 14.560 174.500 14.850 175.665 ;
        RECT 15.450 175.640 15.630 176.310 ;
        RECT 16.375 176.230 18.070 176.400 ;
        RECT 15.800 175.810 16.175 176.140 ;
        RECT 16.345 175.890 17.555 176.060 ;
        RECT 16.345 175.640 16.550 175.890 ;
        RECT 17.725 175.640 18.070 176.230 ;
        RECT 18.245 175.810 18.500 176.370 ;
        RECT 18.670 176.310 19.000 176.845 ;
        RECT 19.215 176.310 19.385 177.050 ;
        RECT 19.595 176.400 19.925 176.870 ;
        RECT 20.095 176.570 20.265 177.050 ;
        RECT 20.435 176.400 20.765 176.870 ;
        RECT 20.935 176.570 21.105 177.050 ;
        RECT 35.590 177.035 39.270 177.205 ;
        RECT 35.735 176.570 35.985 177.035 ;
        RECT 18.670 175.640 18.850 176.310 ;
        RECT 19.595 176.230 21.290 176.400 ;
        RECT 36.155 176.395 36.485 176.865 ;
        RECT 36.655 176.575 36.825 177.035 ;
        RECT 36.995 176.395 37.325 176.865 ;
        RECT 37.495 176.575 37.760 177.035 ;
        RECT 19.020 175.810 19.395 176.140 ;
        RECT 19.565 175.890 20.775 176.060 ;
        RECT 19.565 175.640 19.770 175.890 ;
        RECT 20.945 175.640 21.290 176.230 ;
        RECT 35.720 176.215 37.325 176.395 ;
        RECT 38.220 176.235 38.550 176.865 ;
        RECT 35.720 176.090 35.985 176.215 ;
        RECT 35.640 175.790 35.985 176.090 ;
        RECT 38.220 176.045 38.450 176.235 ;
        RECT 38.720 176.215 38.950 177.035 ;
        RECT 39.450 176.720 41.200 177.240 ;
        RECT 36.155 175.795 38.450 176.045 ;
        RECT 38.620 175.805 38.950 176.045 ;
        RECT 15.090 175.470 16.550 175.640 ;
        RECT 17.215 175.470 18.070 175.640 ;
        RECT 18.310 175.470 19.770 175.640 ;
        RECT 20.435 175.470 21.290 175.640 ;
        RECT 35.720 175.625 35.985 175.790 ;
        RECT 38.220 175.635 38.450 175.795 ;
        RECT 15.090 174.670 15.450 175.470 ;
        RECT 17.215 175.300 17.545 175.470 ;
        RECT 15.995 174.500 16.165 175.300 ;
        RECT 16.375 175.130 17.545 175.300 ;
        RECT 16.375 174.670 16.705 175.130 ;
        RECT 16.875 174.500 17.045 174.960 ;
        RECT 17.215 174.670 17.545 175.130 ;
        RECT 17.715 174.500 17.885 175.300 ;
        RECT 18.310 174.670 18.670 175.470 ;
        RECT 20.435 175.300 20.765 175.470 ;
        RECT 35.720 175.455 37.325 175.625 ;
        RECT 35.720 175.435 36.485 175.455 ;
        RECT 19.215 174.500 19.385 175.300 ;
        RECT 19.595 175.130 20.765 175.300 ;
        RECT 19.595 174.670 19.925 175.130 ;
        RECT 20.095 174.500 20.265 174.960 ;
        RECT 20.435 174.670 20.765 175.130 ;
        RECT 20.935 174.500 21.105 175.300 ;
        RECT 8.035 174.330 21.375 174.500 ;
        RECT 35.775 174.485 35.985 174.945 ;
        RECT 36.155 174.655 36.485 175.435 ;
        RECT 36.655 174.485 36.825 175.285 ;
        RECT 36.995 174.655 37.325 175.455 ;
        RECT 37.495 174.485 37.760 175.625 ;
        RECT 38.220 174.655 38.550 175.635 ;
        RECT 38.720 174.485 38.930 175.625 ;
        RECT 8.130 173.575 8.460 174.330 ;
        RECT 8.640 173.445 8.820 174.160 ;
        RECT 9.025 173.630 9.355 174.330 ;
        RECT 9.565 173.455 9.755 174.160 ;
        RECT 9.925 173.630 10.255 174.330 ;
        RECT 10.425 173.460 10.615 174.160 ;
        RECT 10.785 173.630 11.115 174.330 ;
        RECT 11.350 173.575 11.680 174.330 ;
        RECT 10.425 173.455 11.170 173.460 ;
        RECT 8.160 172.690 8.470 173.310 ;
        RECT 8.640 173.275 9.395 173.445 ;
        RECT 9.185 173.050 9.395 173.275 ;
        RECT 9.565 173.230 11.170 173.455 ;
        RECT 11.860 173.445 12.040 174.160 ;
        RECT 12.245 173.630 12.575 174.330 ;
        RECT 12.785 173.455 12.975 174.160 ;
        RECT 13.145 173.630 13.475 174.330 ;
        RECT 13.645 173.460 13.835 174.160 ;
        RECT 14.005 173.630 14.335 174.330 ;
        RECT 13.645 173.455 14.390 173.460 ;
        RECT 8.640 172.690 9.015 173.020 ;
        RECT 9.185 172.715 10.720 173.050 ;
        RECT 9.185 172.500 9.395 172.715 ;
        RECT 10.890 172.540 11.170 173.230 ;
        RECT 11.380 172.690 11.690 173.310 ;
        RECT 11.860 173.275 12.615 173.445 ;
        RECT 12.405 173.050 12.615 173.275 ;
        RECT 12.785 173.230 14.390 173.455 ;
        RECT 11.860 172.690 12.235 173.020 ;
        RECT 12.405 172.715 13.940 173.050 ;
        RECT 8.130 172.310 9.395 172.500 ;
        RECT 9.565 172.310 11.170 172.540 ;
        RECT 12.405 172.500 12.615 172.715 ;
        RECT 14.110 172.540 14.390 173.230 ;
        RECT 14.560 173.165 14.850 174.330 ;
        RECT 15.090 173.360 15.450 174.160 ;
        RECT 15.995 173.530 16.165 174.330 ;
        RECT 16.375 173.700 16.705 174.160 ;
        RECT 16.875 173.870 17.045 174.330 ;
        RECT 17.215 173.700 17.545 174.160 ;
        RECT 16.375 173.530 17.545 173.700 ;
        RECT 17.715 173.530 17.885 174.330 ;
        RECT 17.215 173.360 17.545 173.530 ;
        RECT 18.310 173.360 18.670 174.160 ;
        RECT 19.215 173.530 19.385 174.330 ;
        RECT 19.595 173.700 19.925 174.160 ;
        RECT 20.095 173.870 20.265 174.330 ;
        RECT 20.435 173.700 20.765 174.160 ;
        RECT 19.595 173.530 20.765 173.700 ;
        RECT 20.935 173.530 21.105 174.330 ;
        RECT 35.590 174.315 39.270 174.485 ;
        RECT 20.435 173.360 20.765 173.530 ;
        RECT 15.090 173.190 16.550 173.360 ;
        RECT 17.215 173.190 18.070 173.360 ;
        RECT 18.310 173.190 19.770 173.360 ;
        RECT 20.435 173.190 21.290 173.360 ;
        RECT 15.025 172.975 15.280 173.020 ;
        RECT 15.015 172.725 15.280 172.975 ;
        RECT 11.350 172.310 12.615 172.500 ;
        RECT 12.785 172.310 14.390 172.540 ;
        RECT 8.130 171.950 8.460 172.310 ;
        RECT 9.565 172.210 9.755 172.310 ;
        RECT 8.990 171.780 9.320 172.140 ;
        RECT 9.925 171.780 10.255 172.140 ;
        RECT 10.425 171.950 10.615 172.310 ;
        RECT 10.785 171.780 11.115 172.140 ;
        RECT 11.350 171.950 11.680 172.310 ;
        RECT 12.785 172.210 12.975 172.310 ;
        RECT 12.210 171.780 12.540 172.140 ;
        RECT 13.145 171.780 13.475 172.140 ;
        RECT 13.645 171.950 13.835 172.310 ;
        RECT 14.005 171.780 14.335 172.140 ;
        RECT 14.560 171.780 14.850 172.505 ;
        RECT 15.025 172.460 15.280 172.725 ;
        RECT 15.450 172.520 15.630 173.190 ;
        RECT 15.800 172.690 16.175 173.020 ;
        RECT 16.345 172.940 16.550 173.190 ;
        RECT 16.345 172.770 17.555 172.940 ;
        RECT 17.725 172.600 18.070 173.190 ;
        RECT 15.040 171.780 15.280 172.290 ;
        RECT 15.450 171.985 15.780 172.520 ;
        RECT 15.995 171.780 16.165 172.520 ;
        RECT 16.375 172.430 18.070 172.600 ;
        RECT 18.245 172.460 18.500 173.020 ;
        RECT 18.670 172.520 18.850 173.190 ;
        RECT 19.020 172.690 19.395 173.020 ;
        RECT 19.565 172.940 19.770 173.190 ;
        RECT 19.565 172.770 20.775 172.940 ;
        RECT 20.945 172.600 21.290 173.190 ;
        RECT 35.685 173.335 36.015 174.145 ;
        RECT 36.185 173.515 36.425 174.315 ;
        RECT 35.685 173.165 36.400 173.335 ;
        RECT 35.680 172.755 36.060 172.995 ;
        RECT 36.230 172.925 36.400 173.165 ;
        RECT 36.605 173.295 36.775 174.145 ;
        RECT 36.945 173.515 37.275 174.315 ;
        RECT 37.445 173.295 37.615 174.145 ;
        RECT 36.605 173.125 37.615 173.295 ;
        RECT 37.785 173.165 38.115 174.315 ;
        RECT 39.450 174.230 39.620 176.720 ;
        RECT 40.160 176.210 40.490 176.380 ;
        RECT 40.020 174.955 40.190 175.995 ;
        RECT 40.460 174.955 40.630 175.995 ;
        RECT 40.160 174.570 40.490 174.740 ;
        RECT 41.030 174.230 41.200 176.720 ;
        RECT 41.600 174.955 41.770 178.995 ;
        RECT 42.040 174.955 42.210 178.995 ;
        RECT 41.740 174.570 42.070 174.740 ;
        RECT 42.610 174.230 42.780 179.720 ;
        RECT 43.320 179.210 43.650 179.380 ;
        RECT 43.180 174.955 43.350 178.995 ;
        RECT 43.620 174.955 43.790 178.995 ;
        RECT 44.190 177.230 44.360 179.720 ;
        RECT 44.900 179.210 45.230 179.380 ;
        RECT 44.760 177.955 44.930 178.995 ;
        RECT 45.200 177.955 45.370 178.995 ;
        RECT 44.900 177.570 45.230 177.740 ;
        RECT 45.770 177.230 45.940 179.720 ;
        RECT 44.190 176.720 45.940 177.230 ;
        RECT 43.320 174.570 43.650 174.740 ;
        RECT 44.190 174.230 44.360 176.720 ;
        RECT 44.900 176.210 45.230 176.380 ;
        RECT 44.760 174.955 44.930 175.995 ;
        RECT 45.200 174.955 45.370 175.995 ;
        RECT 44.900 174.570 45.230 174.740 ;
        RECT 45.770 174.230 45.940 176.720 ;
        RECT 39.450 174.060 45.940 174.230 ;
        RECT 39.455 173.690 45.945 173.700 ;
        RECT 39.340 173.530 46.040 173.690 ;
        RECT 36.230 172.755 36.730 172.925 ;
        RECT 16.375 171.960 16.705 172.430 ;
        RECT 16.875 171.780 17.045 172.260 ;
        RECT 17.215 171.960 17.545 172.430 ;
        RECT 17.715 171.780 17.885 172.260 ;
        RECT 18.260 171.780 18.500 172.290 ;
        RECT 18.670 171.985 19.000 172.520 ;
        RECT 19.215 171.780 19.385 172.520 ;
        RECT 19.595 172.430 21.290 172.600 ;
        RECT 36.230 172.585 36.400 172.755 ;
        RECT 37.120 172.585 37.615 173.125 ;
        RECT 19.595 171.960 19.925 172.430 ;
        RECT 20.095 171.780 20.265 172.260 ;
        RECT 20.435 171.960 20.765 172.430 ;
        RECT 35.765 172.415 36.400 172.585 ;
        RECT 36.605 172.415 37.615 172.585 ;
        RECT 20.935 171.780 21.105 172.260 ;
        RECT 35.765 171.935 35.935 172.415 ;
        RECT 8.035 171.610 21.375 171.780 ;
        RECT 36.115 171.765 36.355 172.245 ;
        RECT 36.605 171.935 36.775 172.415 ;
        RECT 36.945 171.765 37.275 172.245 ;
        RECT 37.445 171.935 37.615 172.415 ;
        RECT 37.785 171.765 38.115 172.565 ;
        RECT 8.130 171.080 8.460 171.440 ;
        RECT 8.990 171.250 9.320 171.610 ;
        RECT 9.925 171.250 10.255 171.610 ;
        RECT 9.565 171.080 9.755 171.180 ;
        RECT 10.425 171.080 10.615 171.440 ;
        RECT 10.785 171.250 11.115 171.610 ;
        RECT 11.350 171.080 11.680 171.440 ;
        RECT 12.210 171.250 12.540 171.610 ;
        RECT 13.145 171.250 13.475 171.610 ;
        RECT 12.785 171.080 12.975 171.180 ;
        RECT 13.645 171.080 13.835 171.440 ;
        RECT 14.005 171.250 14.335 171.610 ;
        RECT 8.130 170.890 9.395 171.080 ;
        RECT 8.215 170.700 8.465 170.715 ;
        RECT 8.160 170.080 8.470 170.700 ;
        RECT 8.640 170.370 9.015 170.700 ;
        RECT 9.185 170.675 9.395 170.890 ;
        RECT 9.565 170.850 11.170 171.080 ;
        RECT 11.350 170.890 12.615 171.080 ;
        RECT 9.185 170.340 10.720 170.675 ;
        RECT 9.185 170.115 9.395 170.340 ;
        RECT 10.890 170.160 11.170 170.850 ;
        RECT 8.640 169.945 9.395 170.115 ;
        RECT 8.130 169.060 8.460 169.815 ;
        RECT 8.640 169.230 8.820 169.945 ;
        RECT 9.565 169.935 11.170 170.160 ;
        RECT 11.380 170.080 11.690 170.700 ;
        RECT 11.860 170.370 12.235 170.700 ;
        RECT 12.405 170.675 12.615 170.890 ;
        RECT 12.785 170.850 14.390 171.080 ;
        RECT 14.560 170.885 14.850 171.610 ;
        RECT 15.040 171.100 15.280 171.610 ;
        RECT 12.405 170.340 13.940 170.675 ;
        RECT 12.405 170.115 12.615 170.340 ;
        RECT 14.110 170.160 14.390 170.850 ;
        RECT 15.025 170.665 15.280 170.930 ;
        RECT 15.015 170.415 15.280 170.665 ;
        RECT 15.025 170.370 15.280 170.415 ;
        RECT 15.450 170.870 15.780 171.405 ;
        RECT 15.995 170.870 16.165 171.610 ;
        RECT 16.375 170.960 16.705 171.430 ;
        RECT 16.875 171.130 17.045 171.610 ;
        RECT 17.215 170.960 17.545 171.430 ;
        RECT 17.715 171.130 17.885 171.610 ;
        RECT 18.260 171.100 18.500 171.610 ;
        RECT 9.025 169.060 9.355 169.760 ;
        RECT 9.565 169.230 9.755 169.935 ;
        RECT 10.425 169.930 11.170 169.935 ;
        RECT 11.860 169.945 12.615 170.115 ;
        RECT 9.925 169.060 10.255 169.760 ;
        RECT 10.425 169.230 10.615 169.930 ;
        RECT 10.785 169.060 11.115 169.760 ;
        RECT 11.350 169.060 11.680 169.815 ;
        RECT 11.860 169.230 12.040 169.945 ;
        RECT 12.785 169.935 14.390 170.160 ;
        RECT 12.245 169.060 12.575 169.760 ;
        RECT 12.785 169.230 12.975 169.935 ;
        RECT 13.645 169.930 14.390 169.935 ;
        RECT 13.145 169.060 13.475 169.760 ;
        RECT 13.645 169.230 13.835 169.930 ;
        RECT 14.005 169.060 14.335 169.760 ;
        RECT 14.560 169.060 14.850 170.225 ;
        RECT 15.450 170.200 15.630 170.870 ;
        RECT 16.375 170.790 18.070 170.960 ;
        RECT 15.800 170.370 16.175 170.700 ;
        RECT 16.345 170.450 17.555 170.620 ;
        RECT 16.345 170.200 16.550 170.450 ;
        RECT 17.725 170.200 18.070 170.790 ;
        RECT 18.245 170.370 18.500 170.930 ;
        RECT 18.670 170.870 19.000 171.405 ;
        RECT 19.215 170.870 19.385 171.610 ;
        RECT 19.595 170.960 19.925 171.430 ;
        RECT 20.095 171.130 20.265 171.610 ;
        RECT 20.435 170.960 20.765 171.430 ;
        RECT 20.935 171.130 21.105 171.610 ;
        RECT 35.590 171.595 38.350 171.765 ;
        RECT 18.670 170.200 18.850 170.870 ;
        RECT 19.595 170.790 21.290 170.960 ;
        RECT 19.020 170.370 19.395 170.700 ;
        RECT 19.565 170.450 20.775 170.620 ;
        RECT 19.565 170.200 19.770 170.450 ;
        RECT 20.945 170.200 21.290 170.790 ;
        RECT 15.090 170.030 16.550 170.200 ;
        RECT 17.215 170.030 18.070 170.200 ;
        RECT 18.310 170.030 19.770 170.200 ;
        RECT 20.435 170.030 21.290 170.200 ;
        RECT 39.340 170.130 39.625 173.530 ;
        RECT 40.165 173.020 40.495 173.190 ;
        RECT 40.025 170.810 40.195 172.850 ;
        RECT 40.465 170.810 40.635 172.850 ;
        RECT 41.035 171.130 41.205 173.530 ;
        RECT 41.745 173.020 42.075 173.190 ;
        RECT 41.605 171.810 41.775 172.850 ;
        RECT 42.045 171.810 42.215 172.850 ;
        RECT 41.745 171.470 42.075 171.640 ;
        RECT 42.615 171.130 42.785 173.530 ;
        RECT 43.325 173.020 43.655 173.190 ;
        RECT 43.185 171.810 43.355 172.850 ;
        RECT 43.625 171.810 43.795 172.850 ;
        RECT 43.325 171.470 43.655 171.640 ;
        RECT 44.195 171.130 44.365 173.530 ;
        RECT 44.905 173.020 45.235 173.190 ;
        RECT 40.165 170.470 40.495 170.640 ;
        RECT 41.035 170.130 44.365 171.130 ;
        RECT 44.765 170.810 44.935 172.850 ;
        RECT 45.205 170.810 45.375 172.850 ;
        RECT 44.905 170.470 45.235 170.640 ;
        RECT 45.775 170.130 46.040 173.530 ;
        RECT 15.090 169.230 15.450 170.030 ;
        RECT 17.215 169.860 17.545 170.030 ;
        RECT 15.995 169.060 16.165 169.860 ;
        RECT 16.375 169.690 17.545 169.860 ;
        RECT 16.375 169.230 16.705 169.690 ;
        RECT 16.875 169.060 17.045 169.520 ;
        RECT 17.215 169.230 17.545 169.690 ;
        RECT 17.715 169.060 17.885 169.860 ;
        RECT 18.310 169.230 18.670 170.030 ;
        RECT 20.435 169.860 20.765 170.030 ;
        RECT 39.340 169.960 46.040 170.130 ;
        RECT 19.215 169.060 19.385 169.860 ;
        RECT 19.595 169.690 20.765 169.860 ;
        RECT 19.595 169.230 19.925 169.690 ;
        RECT 20.095 169.060 20.265 169.520 ;
        RECT 20.435 169.230 20.765 169.690 ;
        RECT 20.935 169.060 21.105 169.860 ;
        RECT 8.035 168.890 21.375 169.060 ;
        RECT 8.130 168.135 8.460 168.890 ;
        RECT 8.640 168.005 8.820 168.720 ;
        RECT 9.025 168.190 9.355 168.890 ;
        RECT 9.565 168.015 9.755 168.720 ;
        RECT 9.925 168.190 10.255 168.890 ;
        RECT 10.425 168.020 10.615 168.720 ;
        RECT 10.785 168.190 11.115 168.890 ;
        RECT 11.350 168.135 11.680 168.890 ;
        RECT 10.425 168.015 11.170 168.020 ;
        RECT 8.160 167.250 8.470 167.870 ;
        RECT 8.640 167.835 9.395 168.005 ;
        RECT 9.185 167.610 9.395 167.835 ;
        RECT 9.565 167.790 11.170 168.015 ;
        RECT 11.860 168.005 12.040 168.720 ;
        RECT 12.245 168.190 12.575 168.890 ;
        RECT 12.785 168.015 12.975 168.720 ;
        RECT 13.145 168.190 13.475 168.890 ;
        RECT 13.645 168.020 13.835 168.720 ;
        RECT 14.005 168.190 14.335 168.890 ;
        RECT 13.645 168.015 14.390 168.020 ;
        RECT 8.640 167.250 9.015 167.580 ;
        RECT 9.185 167.275 10.720 167.610 ;
        RECT 9.185 167.060 9.395 167.275 ;
        RECT 10.890 167.100 11.170 167.790 ;
        RECT 11.380 167.250 11.690 167.870 ;
        RECT 11.860 167.835 12.615 168.005 ;
        RECT 12.405 167.610 12.615 167.835 ;
        RECT 12.785 167.790 14.390 168.015 ;
        RECT 11.860 167.250 12.235 167.580 ;
        RECT 12.405 167.275 13.940 167.610 ;
        RECT 8.130 166.870 9.395 167.060 ;
        RECT 9.565 166.870 11.170 167.100 ;
        RECT 12.405 167.060 12.615 167.275 ;
        RECT 14.110 167.100 14.390 167.790 ;
        RECT 14.560 167.725 14.850 168.890 ;
        RECT 15.090 167.920 15.450 168.720 ;
        RECT 15.995 168.090 16.165 168.890 ;
        RECT 16.375 168.260 16.705 168.720 ;
        RECT 16.875 168.430 17.045 168.890 ;
        RECT 17.215 168.260 17.545 168.720 ;
        RECT 16.375 168.090 17.545 168.260 ;
        RECT 17.715 168.090 17.885 168.890 ;
        RECT 17.215 167.920 17.545 168.090 ;
        RECT 18.310 167.920 18.670 168.720 ;
        RECT 19.215 168.090 19.385 168.890 ;
        RECT 19.595 168.260 19.925 168.720 ;
        RECT 20.095 168.430 20.265 168.890 ;
        RECT 20.435 168.260 20.765 168.720 ;
        RECT 19.595 168.090 20.765 168.260 ;
        RECT 20.935 168.090 21.105 168.890 ;
        RECT 20.435 167.920 20.765 168.090 ;
        RECT 15.090 167.750 16.550 167.920 ;
        RECT 17.215 167.750 18.070 167.920 ;
        RECT 18.310 167.750 19.770 167.920 ;
        RECT 20.435 167.750 21.290 167.920 ;
        RECT 15.025 167.535 15.280 167.580 ;
        RECT 15.015 167.285 15.280 167.535 ;
        RECT 11.350 166.870 12.615 167.060 ;
        RECT 12.785 166.870 14.390 167.100 ;
        RECT 8.130 166.510 8.460 166.870 ;
        RECT 9.565 166.770 9.755 166.870 ;
        RECT 8.990 166.340 9.320 166.700 ;
        RECT 9.925 166.340 10.255 166.700 ;
        RECT 10.425 166.510 10.615 166.870 ;
        RECT 10.785 166.340 11.115 166.700 ;
        RECT 11.350 166.510 11.680 166.870 ;
        RECT 12.785 166.770 12.975 166.870 ;
        RECT 12.210 166.340 12.540 166.700 ;
        RECT 13.145 166.340 13.475 166.700 ;
        RECT 13.645 166.510 13.835 166.870 ;
        RECT 14.005 166.340 14.335 166.700 ;
        RECT 14.560 166.340 14.850 167.065 ;
        RECT 15.025 167.020 15.280 167.285 ;
        RECT 15.450 167.080 15.630 167.750 ;
        RECT 15.800 167.250 16.175 167.580 ;
        RECT 16.345 167.500 16.550 167.750 ;
        RECT 16.345 167.330 17.555 167.500 ;
        RECT 17.725 167.160 18.070 167.750 ;
        RECT 15.040 166.340 15.280 166.850 ;
        RECT 15.450 166.545 15.780 167.080 ;
        RECT 15.995 166.340 16.165 167.080 ;
        RECT 16.375 166.990 18.070 167.160 ;
        RECT 18.245 167.020 18.500 167.580 ;
        RECT 18.670 167.080 18.850 167.750 ;
        RECT 19.020 167.250 19.395 167.580 ;
        RECT 19.565 167.500 19.770 167.750 ;
        RECT 19.565 167.330 20.775 167.500 ;
        RECT 20.945 167.160 21.290 167.750 ;
        RECT 39.340 167.560 40.360 169.960 ;
        RECT 40.920 169.450 41.250 169.620 ;
        RECT 43.020 169.450 43.350 169.620 ;
        RECT 40.760 168.240 40.930 169.280 ;
        RECT 41.240 168.240 41.410 169.280 ;
        RECT 41.810 168.240 41.980 169.280 ;
        RECT 42.290 168.240 42.460 169.280 ;
        RECT 42.860 168.240 43.030 169.280 ;
        RECT 43.340 168.240 43.510 169.280 ;
        RECT 43.910 168.240 44.080 169.280 ;
        RECT 44.390 168.240 44.560 169.280 ;
        RECT 41.970 167.900 42.300 168.070 ;
        RECT 44.070 167.900 44.400 168.070 ;
        RECT 44.960 167.560 46.040 169.960 ;
        RECT 39.340 167.540 46.040 167.560 ;
        RECT 16.375 166.520 16.705 166.990 ;
        RECT 16.875 166.340 17.045 166.820 ;
        RECT 17.215 166.520 17.545 166.990 ;
        RECT 17.715 166.340 17.885 166.820 ;
        RECT 18.260 166.340 18.500 166.850 ;
        RECT 18.670 166.545 19.000 167.080 ;
        RECT 19.215 166.340 19.385 167.080 ;
        RECT 19.595 166.990 21.290 167.160 ;
        RECT 19.595 166.520 19.925 166.990 ;
        RECT 20.095 166.340 20.265 166.820 ;
        RECT 20.435 166.520 20.765 166.990 ;
        RECT 20.935 166.340 21.105 166.820 ;
        RECT 34.640 166.440 46.040 167.540 ;
        RECT 47.420 171.160 48.130 180.770 ;
        RECT 48.610 179.940 50.770 180.290 ;
        RECT 68.610 179.940 70.770 180.290 ;
        RECT 48.610 179.110 50.770 179.460 ;
        RECT 68.610 179.110 70.770 179.460 ;
        RECT 48.610 178.280 50.770 178.630 ;
        RECT 68.610 178.280 70.770 178.630 ;
        RECT 48.610 177.450 50.770 177.800 ;
        RECT 68.610 177.450 70.770 177.800 ;
        RECT 48.610 176.620 50.770 176.970 ;
        RECT 68.610 176.620 70.770 176.970 ;
        RECT 48.610 175.790 50.770 176.140 ;
        RECT 68.610 175.790 70.770 176.140 ;
        RECT 48.610 174.960 50.770 175.310 ;
        RECT 68.610 174.960 70.770 175.310 ;
        RECT 48.610 174.130 50.770 174.480 ;
        RECT 68.610 174.130 70.770 174.480 ;
        RECT 48.610 173.300 50.770 173.650 ;
        RECT 68.610 173.300 70.770 173.650 ;
        RECT 48.610 172.470 50.770 172.820 ;
        RECT 68.610 172.470 70.770 172.820 ;
        RECT 48.610 171.640 50.770 171.990 ;
        RECT 68.610 171.640 70.770 171.990 ;
        RECT 71.250 171.160 71.420 180.770 ;
        RECT 71.780 180.830 102.970 180.940 ;
        RECT 71.780 180.770 73.530 180.830 ;
        RECT 71.780 178.630 71.950 180.770 ;
        RECT 72.350 179.360 72.520 180.400 ;
        RECT 72.790 179.360 72.960 180.400 ;
        RECT 72.490 178.975 72.820 179.145 ;
        RECT 73.360 178.630 73.530 180.770 ;
        RECT 71.780 178.460 73.530 178.630 ;
        RECT 73.890 180.760 102.970 180.830 ;
        RECT 47.420 170.990 71.420 171.160 ;
        RECT 71.780 177.750 73.530 177.920 ;
        RECT 71.780 175.660 71.950 177.750 ;
        RECT 72.490 177.240 72.820 177.410 ;
        RECT 72.350 176.030 72.520 177.070 ;
        RECT 72.790 176.030 72.960 177.070 ;
        RECT 73.360 175.660 73.530 177.750 ;
        RECT 71.780 175.490 73.530 175.660 ;
        RECT 47.420 169.660 48.070 170.990 ;
        RECT 54.870 169.750 60.970 170.180 ;
        RECT 47.420 169.490 54.250 169.660 ;
        RECT 8.035 166.170 21.375 166.340 ;
        RECT 47.420 166.090 48.130 169.490 ;
        RECT 48.690 168.980 49.020 169.150 ;
        RECT 49.650 168.980 49.980 169.150 ;
        RECT 48.530 166.770 48.700 168.810 ;
        RECT 49.010 166.770 49.180 168.810 ;
        RECT 49.490 166.770 49.660 168.810 ;
        RECT 49.970 166.770 50.140 168.810 ;
        RECT 50.450 166.770 50.620 168.810 ;
        RECT 49.170 166.430 49.500 166.600 ;
        RECT 50.130 166.430 50.460 166.600 ;
        RECT 51.020 166.090 51.190 169.490 ;
        RECT 51.750 168.980 52.080 169.150 ;
        RECT 52.710 168.980 53.040 169.150 ;
        RECT 51.590 166.770 51.760 168.810 ;
        RECT 52.070 166.770 52.240 168.810 ;
        RECT 52.550 166.770 52.720 168.810 ;
        RECT 53.030 166.770 53.200 168.810 ;
        RECT 53.510 166.770 53.680 168.810 ;
        RECT 52.230 166.430 52.560 166.600 ;
        RECT 53.190 166.430 53.520 166.600 ;
        RECT 54.080 166.090 54.250 169.490 ;
        RECT 47.420 165.920 54.250 166.090 ;
        RECT 54.770 169.580 61.060 169.750 ;
        RECT 54.770 166.090 54.940 169.580 ;
        RECT 55.500 169.070 55.830 169.240 ;
        RECT 56.460 169.070 56.790 169.240 ;
        RECT 55.340 166.815 55.510 168.855 ;
        RECT 55.820 166.815 55.990 168.855 ;
        RECT 56.300 166.815 56.470 168.855 ;
        RECT 56.780 166.815 56.950 168.855 ;
        RECT 57.260 166.815 57.430 168.855 ;
        RECT 55.980 166.430 56.310 166.600 ;
        RECT 56.940 166.430 57.270 166.600 ;
        RECT 57.830 166.090 58.000 169.580 ;
        RECT 58.560 169.070 58.890 169.240 ;
        RECT 59.520 169.070 59.850 169.240 ;
        RECT 58.400 166.815 58.570 168.855 ;
        RECT 58.880 166.815 59.050 168.855 ;
        RECT 59.360 166.815 59.530 168.855 ;
        RECT 59.840 166.815 60.010 168.855 ;
        RECT 60.320 166.815 60.490 168.855 ;
        RECT 59.040 166.430 59.370 166.600 ;
        RECT 60.000 166.430 60.330 166.600 ;
        RECT 60.890 166.090 61.060 169.580 ;
        RECT 54.770 165.920 61.060 166.090 ;
        RECT 63.060 169.390 66.290 169.560 ;
        RECT 63.060 166.090 63.230 169.390 ;
        RECT 63.790 168.880 64.120 169.050 ;
        RECT 64.750 168.880 65.080 169.050 ;
        RECT 63.630 166.770 63.800 168.710 ;
        RECT 64.110 166.770 64.280 168.710 ;
        RECT 64.590 166.770 64.760 168.710 ;
        RECT 65.070 166.770 65.240 168.710 ;
        RECT 65.550 166.770 65.720 168.710 ;
        RECT 64.270 166.430 64.600 166.600 ;
        RECT 65.230 166.430 65.560 166.600 ;
        RECT 66.120 166.090 66.290 169.390 ;
        RECT 63.060 165.980 66.290 166.090 ;
        RECT 68.330 168.100 71.420 168.270 ;
        RECT 68.330 166.150 68.500 168.100 ;
        RECT 69.000 167.010 69.170 167.550 ;
        RECT 69.790 167.010 69.960 167.550 ;
        RECT 70.580 167.010 70.750 167.550 ;
        RECT 69.230 166.670 69.730 166.840 ;
        RECT 70.020 166.670 70.520 166.840 ;
        RECT 71.250 166.150 71.420 168.100 ;
        RECT 68.330 165.980 71.420 166.150 ;
        RECT 71.780 166.090 71.950 175.490 ;
        RECT 72.490 174.980 72.820 175.150 ;
        RECT 72.350 166.770 72.520 174.810 ;
        RECT 72.790 167.130 72.960 174.810 ;
        RECT 73.360 167.130 73.530 175.490 ;
        RECT 72.790 166.830 73.530 167.130 ;
        RECT 72.790 166.770 72.960 166.830 ;
        RECT 72.490 166.430 72.820 166.600 ;
        RECT 73.220 166.090 73.530 166.830 ;
        RECT 71.780 165.980 73.530 166.090 ;
        RECT 63.060 165.920 73.530 165.980 ;
        RECT 73.890 166.090 74.060 180.760 ;
        RECT 75.115 180.250 75.445 180.420 ;
        RECT 76.095 180.250 76.425 180.420 ;
        RECT 77.075 180.250 77.405 180.420 ;
        RECT 78.055 180.250 78.385 180.420 ;
        RECT 74.460 173.995 74.630 180.035 ;
        RECT 74.950 173.995 75.120 180.035 ;
        RECT 75.440 173.995 75.610 180.035 ;
        RECT 75.930 173.995 76.100 180.035 ;
        RECT 76.420 173.995 76.590 180.035 ;
        RECT 76.910 173.995 77.080 180.035 ;
        RECT 77.400 173.995 77.570 180.035 ;
        RECT 77.890 173.995 78.060 180.035 ;
        RECT 78.380 173.995 78.550 180.035 ;
        RECT 74.625 173.610 74.955 173.780 ;
        RECT 75.605 173.610 75.935 173.780 ;
        RECT 76.585 173.610 76.915 173.780 ;
        RECT 77.565 173.610 77.895 173.780 ;
        RECT 74.625 173.070 74.955 173.240 ;
        RECT 75.605 173.070 75.935 173.240 ;
        RECT 76.585 173.070 76.915 173.240 ;
        RECT 77.565 173.070 77.895 173.240 ;
        RECT 74.460 166.815 74.630 172.855 ;
        RECT 74.950 166.815 75.120 172.855 ;
        RECT 75.440 166.815 75.610 172.855 ;
        RECT 75.930 166.815 76.100 172.855 ;
        RECT 76.420 166.815 76.590 172.855 ;
        RECT 76.910 166.815 77.080 172.855 ;
        RECT 77.400 166.815 77.570 172.855 ;
        RECT 77.890 166.815 78.060 172.855 ;
        RECT 78.380 166.815 78.550 172.855 ;
        RECT 75.115 166.430 75.445 166.600 ;
        RECT 76.095 166.430 76.425 166.600 ;
        RECT 77.075 166.430 77.405 166.600 ;
        RECT 78.055 166.430 78.385 166.600 ;
        RECT 78.950 166.090 79.120 180.760 ;
        RECT 80.175 180.250 80.505 180.420 ;
        RECT 81.155 180.250 81.485 180.420 ;
        RECT 82.135 180.250 82.465 180.420 ;
        RECT 83.115 180.250 83.445 180.420 ;
        RECT 79.520 173.995 79.690 180.035 ;
        RECT 80.010 173.995 80.180 180.035 ;
        RECT 80.500 173.995 80.670 180.035 ;
        RECT 80.990 173.995 81.160 180.035 ;
        RECT 81.480 173.995 81.650 180.035 ;
        RECT 81.970 173.995 82.140 180.035 ;
        RECT 82.460 173.995 82.630 180.035 ;
        RECT 82.950 173.995 83.120 180.035 ;
        RECT 83.440 173.995 83.610 180.035 ;
        RECT 79.685 173.610 80.015 173.780 ;
        RECT 80.665 173.610 80.995 173.780 ;
        RECT 81.645 173.610 81.975 173.780 ;
        RECT 82.625 173.610 82.955 173.780 ;
        RECT 79.685 173.070 80.015 173.240 ;
        RECT 80.665 173.070 80.995 173.240 ;
        RECT 81.645 173.070 81.975 173.240 ;
        RECT 82.625 173.070 82.955 173.240 ;
        RECT 79.520 166.815 79.690 172.855 ;
        RECT 80.010 166.815 80.180 172.855 ;
        RECT 80.500 166.815 80.670 172.855 ;
        RECT 80.990 166.815 81.160 172.855 ;
        RECT 81.480 166.815 81.650 172.855 ;
        RECT 81.970 166.815 82.140 172.855 ;
        RECT 82.460 166.815 82.630 172.855 ;
        RECT 82.950 166.815 83.120 172.855 ;
        RECT 83.440 166.815 83.610 172.855 ;
        RECT 84.000 171.270 84.180 180.760 ;
        RECT 84.800 180.250 85.300 180.420 ;
        RECT 86.160 180.250 86.660 180.420 ;
        RECT 87.520 180.250 88.020 180.420 ;
        RECT 88.880 180.250 89.380 180.420 ;
        RECT 90.240 180.250 90.740 180.420 ;
        RECT 91.600 180.250 92.100 180.420 ;
        RECT 92.960 180.250 93.460 180.420 ;
        RECT 94.320 180.250 94.820 180.420 ;
        RECT 95.680 180.250 96.180 180.420 ;
        RECT 97.040 180.250 97.540 180.420 ;
        RECT 98.400 180.250 98.900 180.420 ;
        RECT 99.760 180.250 100.260 180.420 ;
        RECT 101.120 180.250 101.620 180.420 ;
        RECT 84.570 171.995 84.740 180.035 ;
        RECT 85.360 171.995 85.530 180.035 ;
        RECT 85.930 171.995 86.100 180.035 ;
        RECT 86.720 171.995 86.890 180.035 ;
        RECT 87.290 171.995 87.460 180.035 ;
        RECT 88.080 171.995 88.250 180.035 ;
        RECT 88.650 171.995 88.820 180.035 ;
        RECT 89.440 171.995 89.610 180.035 ;
        RECT 90.010 171.995 90.180 180.035 ;
        RECT 90.800 171.995 90.970 180.035 ;
        RECT 91.370 171.995 91.540 180.035 ;
        RECT 92.160 171.995 92.330 180.035 ;
        RECT 92.730 171.995 92.900 180.035 ;
        RECT 93.520 171.995 93.690 180.035 ;
        RECT 94.090 171.995 94.260 180.035 ;
        RECT 94.880 171.995 95.050 180.035 ;
        RECT 95.450 171.995 95.620 180.035 ;
        RECT 96.240 171.995 96.410 180.035 ;
        RECT 96.810 171.995 96.980 180.035 ;
        RECT 97.600 171.995 97.770 180.035 ;
        RECT 98.170 171.995 98.340 180.035 ;
        RECT 98.960 171.995 99.130 180.035 ;
        RECT 99.530 171.995 99.700 180.035 ;
        RECT 100.320 171.995 100.490 180.035 ;
        RECT 100.890 171.995 101.060 180.035 ;
        RECT 101.680 171.995 101.850 180.035 ;
        RECT 84.800 171.610 85.300 171.780 ;
        RECT 86.160 171.610 86.660 171.780 ;
        RECT 87.520 171.610 88.020 171.780 ;
        RECT 88.880 171.610 89.380 171.780 ;
        RECT 90.240 171.610 90.740 171.780 ;
        RECT 91.600 171.610 92.100 171.780 ;
        RECT 92.960 171.610 93.460 171.780 ;
        RECT 94.320 171.610 94.820 171.780 ;
        RECT 95.680 171.610 96.180 171.780 ;
        RECT 97.040 171.610 97.540 171.780 ;
        RECT 98.400 171.610 98.900 171.780 ;
        RECT 99.760 171.610 100.260 171.780 ;
        RECT 101.120 171.610 101.620 171.780 ;
        RECT 102.250 171.270 102.970 180.760 ;
        RECT 84.000 171.100 102.970 171.270 ;
        RECT 80.175 166.430 80.505 166.600 ;
        RECT 81.155 166.430 81.485 166.600 ;
        RECT 82.135 166.430 82.465 166.600 ;
        RECT 83.115 166.430 83.445 166.600 ;
        RECT 84.010 166.090 84.180 171.100 ;
        RECT 84.670 170.450 90.660 170.620 ;
        RECT 84.670 167.050 84.840 170.450 ;
        RECT 86.450 169.940 86.780 170.110 ;
        RECT 88.550 169.940 88.880 170.110 ;
        RECT 85.240 167.730 85.410 169.770 ;
        RECT 85.720 167.730 85.890 169.770 ;
        RECT 86.290 167.730 86.460 169.770 ;
        RECT 86.770 167.730 86.940 169.770 ;
        RECT 87.340 167.730 87.510 169.770 ;
        RECT 87.820 167.730 87.990 169.770 ;
        RECT 88.390 167.730 88.560 169.770 ;
        RECT 88.870 167.730 89.040 169.770 ;
        RECT 89.440 167.730 89.610 169.770 ;
        RECT 89.920 167.730 90.090 169.770 ;
        RECT 85.400 167.390 85.730 167.560 ;
        RECT 87.500 167.390 87.830 167.560 ;
        RECT 89.600 167.390 89.930 167.560 ;
        RECT 90.490 167.050 90.660 170.450 ;
        RECT 91.910 168.960 92.080 171.100 ;
        RECT 92.480 169.690 92.650 170.730 ;
        RECT 93.770 169.690 93.940 170.730 ;
        RECT 95.060 169.690 95.230 170.730 ;
        RECT 95.630 170.685 102.970 171.100 ;
        RECT 95.630 170.680 101.270 170.685 ;
        RECT 92.710 169.305 93.710 169.475 ;
        RECT 94.000 169.305 95.000 169.475 ;
        RECT 95.630 168.960 95.800 170.680 ;
        RECT 91.910 168.790 95.800 168.960 ;
        RECT 101.370 169.535 101.700 170.515 ;
        RECT 101.870 169.545 102.080 170.685 ;
        RECT 102.320 170.530 102.970 170.685 ;
        RECT 109.245 173.525 109.745 185.015 ;
        RECT 141.435 184.715 141.605 185.015 ;
        RECT 141.815 184.815 144.575 184.985 ;
        RECT 110.225 184.505 120.225 184.675 ;
        RECT 120.515 184.505 130.515 184.675 ;
        RECT 130.805 184.505 140.805 184.675 ;
        RECT 109.995 174.250 110.165 184.290 ;
        RECT 120.285 174.250 120.455 184.290 ;
        RECT 130.575 174.250 130.745 184.290 ;
        RECT 140.865 174.250 141.035 184.290 ;
        RECT 110.225 173.865 120.225 174.035 ;
        RECT 120.515 173.865 130.515 174.035 ;
        RECT 130.805 173.865 140.805 174.035 ;
        RECT 141.395 173.525 141.605 184.715 ;
        RECT 142.145 184.015 142.475 184.645 ;
        RECT 142.145 183.415 142.375 184.015 ;
        RECT 142.645 183.995 142.875 184.815 ;
        RECT 143.280 184.015 143.975 184.645 ;
        RECT 144.180 184.015 144.490 184.815 ;
        RECT 142.545 183.585 142.875 183.825 ;
        RECT 143.300 183.575 143.635 183.825 ;
        RECT 143.805 183.415 143.975 184.015 ;
        RECT 144.145 183.575 144.480 183.845 ;
        RECT 142.145 182.435 142.475 183.415 ;
        RECT 142.645 182.265 142.855 183.405 ;
        RECT 143.280 182.265 143.540 183.405 ;
        RECT 143.710 182.435 144.040 183.415 ;
        RECT 144.210 182.265 144.490 183.405 ;
        RECT 141.815 182.095 144.575 182.265 ;
        RECT 142.145 180.945 142.475 181.925 ;
        RECT 142.645 180.955 142.855 182.095 ;
        RECT 143.280 180.955 143.540 182.095 ;
        RECT 143.710 180.945 144.040 181.925 ;
        RECT 144.210 180.955 144.490 182.095 ;
        RECT 142.145 180.345 142.375 180.945 ;
        RECT 142.555 180.775 142.860 180.780 ;
        RECT 142.545 180.535 142.875 180.775 ;
        RECT 143.300 180.535 143.635 180.785 ;
        RECT 142.145 179.715 142.475 180.345 ;
        RECT 142.645 179.545 142.875 180.365 ;
        RECT 143.805 180.345 143.975 180.945 ;
        RECT 144.145 180.515 144.480 180.785 ;
        RECT 143.280 179.715 143.975 180.345 ;
        RECT 144.180 179.545 144.490 180.345 ;
        RECT 141.815 179.375 145.035 179.545 ;
        RECT 142.145 178.575 142.475 179.205 ;
        RECT 142.145 177.975 142.375 178.575 ;
        RECT 142.645 178.555 142.875 179.375 ;
        RECT 143.290 178.865 144.520 179.205 ;
        RECT 144.690 178.885 144.945 179.375 ;
        RECT 143.290 178.635 143.620 178.865 ;
        RECT 142.545 178.145 142.875 178.385 ;
        RECT 143.280 178.135 143.595 178.465 ;
        RECT 143.795 178.135 144.170 178.695 ;
        RECT 142.145 176.995 142.475 177.975 ;
        RECT 144.340 177.965 144.520 178.865 ;
        RECT 144.705 178.515 144.925 178.715 ;
        RECT 144.705 178.165 145.045 178.515 ;
        RECT 144.705 178.135 144.925 178.165 ;
        RECT 142.645 176.825 142.855 177.965 ;
        RECT 143.290 177.795 144.520 177.965 ;
        RECT 143.290 176.995 143.620 177.795 ;
        RECT 143.790 176.825 144.020 177.625 ;
        RECT 144.190 176.995 144.520 177.795 ;
        RECT 144.690 176.825 144.945 177.965 ;
        RECT 141.815 176.655 145.035 176.825 ;
        RECT 142.155 175.515 142.365 176.655 ;
        RECT 142.535 176.060 142.865 176.485 ;
        RECT 142.535 175.820 142.870 176.060 ;
        RECT 142.535 175.505 142.865 175.820 ;
        RECT 143.535 175.515 143.745 176.655 ;
        RECT 143.915 175.505 144.245 176.485 ;
        RECT 142.135 175.095 142.465 175.335 ;
        RECT 142.135 174.105 142.365 174.925 ;
        RECT 142.635 174.905 142.865 175.505 ;
        RECT 143.515 175.095 143.845 175.335 ;
        RECT 142.535 174.275 142.865 174.905 ;
        RECT 143.515 174.105 143.745 174.925 ;
        RECT 144.015 174.905 144.245 175.505 ;
        RECT 143.915 174.275 144.245 174.905 ;
        RECT 141.815 173.935 144.575 174.105 ;
        RECT 109.245 173.355 141.605 173.525 ;
        RECT 101.370 168.935 101.600 169.535 ;
        RECT 101.770 169.125 102.100 169.365 ;
        RECT 101.370 168.305 101.700 168.935 ;
        RECT 101.870 168.135 102.100 168.955 ;
        RECT 101.040 168.080 102.420 168.135 ;
        RECT 101.040 167.965 102.970 168.080 ;
        RECT 84.670 166.880 90.660 167.050 ;
        RECT 73.890 165.920 84.180 166.090 ;
        RECT 84.720 165.980 90.620 166.880 ;
        RECT 101.070 165.980 102.970 167.965 ;
        RECT 47.420 165.580 54.220 165.920 ;
        RECT 63.120 165.580 73.520 165.920 ;
        RECT 84.720 165.580 102.970 165.980 ;
        RECT 47.420 164.880 102.970 165.580 ;
        RECT 109.245 161.865 109.745 173.355 ;
        RECT 110.225 172.845 120.225 173.015 ;
        RECT 120.515 172.845 130.515 173.015 ;
        RECT 130.805 172.845 140.805 173.015 ;
        RECT 141.395 172.655 141.605 173.355 ;
        RECT 109.995 162.590 110.165 172.630 ;
        RECT 120.285 162.590 120.455 172.630 ;
        RECT 130.575 162.590 130.745 172.630 ;
        RECT 140.865 162.590 141.035 172.630 ;
        RECT 141.395 172.485 144.665 172.655 ;
        RECT 141.395 170.575 141.605 172.485 ;
        RECT 142.645 171.975 142.975 172.145 ;
        RECT 143.605 171.975 143.935 172.145 ;
        RECT 142.005 171.300 142.175 171.760 ;
        RECT 142.485 171.300 142.655 171.760 ;
        RECT 142.965 171.300 143.135 171.760 ;
        RECT 143.445 171.300 143.615 171.760 ;
        RECT 143.925 171.300 144.095 171.760 ;
        RECT 142.165 170.915 142.495 171.085 ;
        RECT 143.125 170.915 143.455 171.085 ;
        RECT 144.495 170.575 144.665 172.485 ;
        RECT 141.395 170.405 144.665 170.575 ;
        RECT 141.395 168.495 141.605 170.405 ;
        RECT 142.165 169.895 142.495 170.065 ;
        RECT 143.125 169.895 143.455 170.065 ;
        RECT 142.005 169.220 142.175 169.680 ;
        RECT 142.485 169.220 142.655 169.680 ;
        RECT 142.965 169.220 143.135 169.680 ;
        RECT 143.445 169.220 143.615 169.680 ;
        RECT 143.925 169.220 144.095 169.680 ;
        RECT 142.645 168.835 142.975 169.005 ;
        RECT 143.605 168.835 143.935 169.005 ;
        RECT 144.495 168.495 144.665 170.405 ;
        RECT 141.395 168.325 144.665 168.495 ;
        RECT 141.395 168.315 141.605 168.325 ;
        RECT 110.225 162.205 120.225 162.375 ;
        RECT 120.515 162.205 130.515 162.375 ;
        RECT 130.805 162.205 140.805 162.375 ;
        RECT 141.435 161.865 141.605 168.315 ;
        RECT 141.995 167.005 142.445 167.165 ;
        RECT 141.975 166.835 144.725 167.005 ;
        RECT 141.975 165.015 142.145 166.835 ;
        RECT 142.705 166.325 143.035 166.495 ;
        RECT 143.665 166.325 143.995 166.495 ;
        RECT 142.545 165.695 142.715 166.155 ;
        RECT 143.025 165.695 143.195 166.155 ;
        RECT 143.505 165.695 143.675 166.155 ;
        RECT 143.985 165.695 144.155 166.155 ;
        RECT 143.185 165.355 143.515 165.525 ;
        RECT 144.555 165.015 144.725 166.835 ;
        RECT 141.975 164.845 144.725 165.015 ;
        RECT 141.975 163.025 142.145 164.845 ;
        RECT 143.185 164.335 143.515 164.505 ;
        RECT 142.545 163.705 142.715 164.165 ;
        RECT 143.025 163.705 143.195 164.165 ;
        RECT 143.505 163.705 143.675 164.165 ;
        RECT 143.985 163.705 144.155 164.165 ;
        RECT 142.705 163.365 143.035 163.535 ;
        RECT 143.665 163.365 143.995 163.535 ;
        RECT 144.555 163.025 144.725 164.845 ;
        RECT 141.975 162.855 144.725 163.025 ;
        RECT 109.245 161.695 141.605 161.865 ;
        RECT 109.245 161.515 141.445 161.695 ;
        RECT 20.470 160.035 23.970 160.150 ;
        RECT 137.145 160.035 140.645 160.150 ;
        RECT 20.470 160.030 24.000 160.035 ;
        RECT 137.115 160.030 140.645 160.035 ;
        RECT 20.205 159.860 37.475 160.030 ;
        RECT 20.350 159.395 20.600 159.860 ;
        RECT 20.770 159.220 21.100 159.690 ;
        RECT 21.270 159.400 21.440 159.860 ;
        RECT 21.610 159.220 21.940 159.690 ;
        RECT 22.110 159.400 22.375 159.860 ;
        RECT 20.335 159.040 21.940 159.220 ;
        RECT 22.650 159.040 22.860 159.860 ;
        RECT 23.030 159.060 23.360 159.690 ;
        RECT 20.335 158.450 20.600 159.040 ;
        RECT 23.030 158.870 23.280 159.060 ;
        RECT 23.530 159.040 23.760 159.860 ;
        RECT 24.255 159.830 37.475 159.860 ;
        RECT 20.770 158.620 23.280 158.870 ;
        RECT 23.450 158.840 23.780 158.870 ;
        RECT 23.450 158.670 24.005 158.840 ;
        RECT 23.450 158.620 23.780 158.670 ;
        RECT 23.030 158.460 23.280 158.620 ;
        RECT 20.335 158.280 21.940 158.450 ;
        RECT 20.335 158.260 21.100 158.280 ;
        RECT 20.390 157.310 20.600 157.770 ;
        RECT 20.770 157.480 21.100 158.260 ;
        RECT 21.270 157.310 21.440 158.110 ;
        RECT 21.610 157.480 21.940 158.280 ;
        RECT 22.110 157.310 22.375 158.450 ;
        RECT 22.650 157.310 22.860 158.450 ;
        RECT 23.030 157.480 23.360 158.460 ;
        RECT 23.530 157.310 23.760 158.450 ;
        RECT 20.205 157.140 23.885 157.310 ;
        RECT 20.590 155.975 21.235 157.140 ;
        RECT 21.715 156.000 21.980 157.140 ;
        RECT 22.150 156.170 22.480 156.970 ;
        RECT 22.650 156.340 22.820 157.140 ;
        RECT 22.990 156.190 23.320 156.970 ;
        RECT 23.490 156.680 23.700 157.140 ;
        RECT 22.990 156.170 23.755 156.190 ;
        RECT 22.150 156.000 23.755 156.170 ;
        RECT 21.690 155.580 23.320 155.830 ;
        RECT 23.490 155.410 23.755 156.000 ;
        RECT 22.150 155.230 23.755 155.410 ;
        RECT 21.715 154.590 21.980 155.050 ;
        RECT 22.150 154.760 22.480 155.230 ;
        RECT 22.650 154.590 22.820 155.050 ;
        RECT 22.990 154.760 23.320 155.230 ;
        RECT 23.490 154.590 23.740 155.055 ;
        RECT 21.585 154.460 23.885 154.590 ;
        RECT 24.255 154.460 24.425 159.830 ;
        RECT 24.825 155.140 24.995 159.180 ;
        RECT 25.305 155.140 25.475 159.180 ;
        RECT 25.785 155.140 25.955 159.180 ;
        RECT 24.985 154.800 25.315 154.970 ;
        RECT 26.355 154.460 26.525 159.830 ;
        RECT 27.085 159.350 27.415 159.520 ;
        RECT 26.925 155.140 27.095 159.180 ;
        RECT 27.405 155.140 27.575 159.180 ;
        RECT 27.885 155.140 28.055 159.180 ;
        RECT 28.455 154.460 28.625 159.830 ;
        RECT 29.025 155.140 29.195 159.180 ;
        RECT 29.505 155.140 29.675 159.180 ;
        RECT 29.985 155.140 30.155 159.180 ;
        RECT 29.185 154.800 29.515 154.970 ;
        RECT 30.555 154.460 30.725 159.830 ;
        RECT 21.585 154.420 23.890 154.460 ;
        RECT 21.700 154.290 23.890 154.420 ;
        RECT 24.255 154.290 30.725 154.460 ;
        RECT 31.055 154.100 31.225 159.830 ;
        RECT 31.955 159.170 32.855 159.340 ;
        RECT 31.725 154.960 31.895 159.000 ;
        RECT 32.915 154.960 33.085 159.000 ;
        RECT 31.955 154.620 32.855 154.790 ;
        RECT 33.585 154.100 33.755 159.830 ;
        RECT 34.485 159.170 35.385 159.340 ;
        RECT 35.675 159.170 36.575 159.340 ;
        RECT 34.255 154.960 34.425 159.000 ;
        RECT 35.445 154.960 35.615 159.000 ;
        RECT 36.635 154.960 36.805 159.000 ;
        RECT 34.485 154.620 35.385 154.790 ;
        RECT 35.675 154.620 36.575 154.790 ;
        RECT 37.305 154.100 37.475 159.830 ;
        RECT 37.895 159.860 74.425 160.030 ;
        RECT 37.895 159.095 38.065 159.860 ;
        RECT 37.895 155.700 38.070 159.095 ;
        RECT 37.895 154.370 38.065 155.700 ;
        RECT 38.465 155.095 38.635 159.135 ;
        RECT 38.945 155.095 39.115 159.135 ;
        RECT 39.425 155.095 39.595 159.135 ;
        RECT 39.905 155.095 40.075 159.135 ;
        RECT 40.385 155.095 40.555 159.135 ;
        RECT 40.955 157.370 41.125 159.860 ;
        RECT 41.665 159.350 41.995 159.520 ;
        RECT 41.525 158.095 41.695 159.135 ;
        RECT 41.965 158.095 42.135 159.135 ;
        RECT 42.535 157.370 42.705 159.860 ;
        RECT 43.335 159.350 58.335 159.520 ;
        RECT 58.625 159.350 73.625 159.520 ;
        RECT 40.955 157.200 42.705 157.370 ;
        RECT 38.625 154.710 38.955 154.880 ;
        RECT 39.585 154.710 39.915 154.880 ;
        RECT 40.955 154.370 41.125 157.200 ;
        RECT 37.895 154.200 41.125 154.370 ;
        RECT 38.335 154.100 40.335 154.200 ;
        RECT 31.055 153.930 37.475 154.100 ;
        RECT 42.535 149.690 42.705 157.200 ;
        RECT 43.105 155.345 43.275 159.135 ;
        RECT 58.395 155.345 58.565 159.135 ;
        RECT 73.685 155.345 73.855 159.135 ;
        RECT 74.255 159.125 74.425 159.860 ;
        RECT 86.690 159.860 123.220 160.030 ;
        RECT 86.690 159.125 86.860 159.860 ;
        RECT 87.490 159.350 102.490 159.520 ;
        RECT 102.780 159.350 117.780 159.520 ;
        RECT 74.255 155.730 74.430 159.125 ;
        RECT 86.685 155.730 86.860 159.125 ;
        RECT 43.335 154.960 58.335 155.130 ;
        RECT 58.625 154.960 73.625 155.130 ;
        RECT 43.335 154.420 58.335 154.590 ;
        RECT 58.625 154.420 73.625 154.590 ;
        RECT 43.105 150.415 43.275 154.205 ;
        RECT 58.395 150.415 58.565 154.205 ;
        RECT 73.685 150.415 73.855 154.205 ;
        RECT 43.335 150.030 58.335 150.200 ;
        RECT 58.625 150.030 73.625 150.200 ;
        RECT 43.505 149.690 58.340 149.715 ;
        RECT 74.255 149.690 74.425 155.730 ;
        RECT 42.535 149.520 74.425 149.690 ;
        RECT 86.690 149.690 86.860 155.730 ;
        RECT 87.260 155.345 87.430 159.135 ;
        RECT 102.550 155.345 102.720 159.135 ;
        RECT 117.840 155.345 118.010 159.135 ;
        RECT 118.410 157.370 118.580 159.860 ;
        RECT 119.120 159.350 119.450 159.520 ;
        RECT 118.980 158.095 119.150 159.135 ;
        RECT 119.420 158.095 119.590 159.135 ;
        RECT 119.990 157.370 120.160 159.860 ;
        RECT 118.410 157.200 120.160 157.370 ;
        RECT 87.490 154.960 102.490 155.130 ;
        RECT 102.780 154.960 117.780 155.130 ;
        RECT 87.490 154.420 102.490 154.590 ;
        RECT 102.780 154.420 117.780 154.590 ;
        RECT 87.260 150.415 87.430 154.205 ;
        RECT 102.550 150.415 102.720 154.205 ;
        RECT 117.840 150.415 118.010 154.205 ;
        RECT 87.490 150.030 102.490 150.200 ;
        RECT 102.780 150.030 117.780 150.200 ;
        RECT 102.775 149.690 117.610 149.715 ;
        RECT 118.410 149.690 118.580 157.200 ;
        RECT 119.990 154.370 120.160 157.200 ;
        RECT 120.560 155.095 120.730 159.135 ;
        RECT 121.040 155.095 121.210 159.135 ;
        RECT 121.520 155.095 121.690 159.135 ;
        RECT 122.000 155.095 122.170 159.135 ;
        RECT 122.480 155.095 122.650 159.135 ;
        RECT 123.050 159.095 123.220 159.860 ;
        RECT 123.045 155.700 123.220 159.095 ;
        RECT 121.200 154.710 121.530 154.880 ;
        RECT 122.160 154.710 122.490 154.880 ;
        RECT 123.050 154.370 123.220 155.700 ;
        RECT 119.990 154.200 123.220 154.370 ;
        RECT 123.640 159.860 140.910 160.030 ;
        RECT 123.640 159.830 136.860 159.860 ;
        RECT 120.780 154.100 122.780 154.200 ;
        RECT 123.640 154.100 123.810 159.830 ;
        RECT 124.540 159.170 125.440 159.340 ;
        RECT 125.730 159.170 126.630 159.340 ;
        RECT 124.310 154.960 124.480 159.000 ;
        RECT 125.500 154.960 125.670 159.000 ;
        RECT 126.690 154.960 126.860 159.000 ;
        RECT 124.540 154.620 125.440 154.790 ;
        RECT 125.730 154.620 126.630 154.790 ;
        RECT 127.360 154.100 127.530 159.830 ;
        RECT 128.260 159.170 129.160 159.340 ;
        RECT 128.030 154.960 128.200 159.000 ;
        RECT 129.220 154.960 129.390 159.000 ;
        RECT 128.260 154.620 129.160 154.790 ;
        RECT 129.890 154.100 130.060 159.830 ;
        RECT 130.390 154.460 130.560 159.830 ;
        RECT 130.960 155.140 131.130 159.180 ;
        RECT 131.440 155.140 131.610 159.180 ;
        RECT 131.920 155.140 132.090 159.180 ;
        RECT 131.600 154.800 131.930 154.970 ;
        RECT 132.490 154.460 132.660 159.830 ;
        RECT 133.700 159.350 134.030 159.520 ;
        RECT 133.060 155.140 133.230 159.180 ;
        RECT 133.540 155.140 133.710 159.180 ;
        RECT 134.020 155.140 134.190 159.180 ;
        RECT 134.590 154.460 134.760 159.830 ;
        RECT 135.160 155.140 135.330 159.180 ;
        RECT 135.640 155.140 135.810 159.180 ;
        RECT 136.120 155.140 136.290 159.180 ;
        RECT 135.800 154.800 136.130 154.970 ;
        RECT 136.690 154.460 136.860 159.830 ;
        RECT 137.355 159.040 137.585 159.860 ;
        RECT 137.755 159.060 138.085 159.690 ;
        RECT 137.835 158.870 138.085 159.060 ;
        RECT 138.255 159.040 138.465 159.860 ;
        RECT 138.740 159.400 139.005 159.860 ;
        RECT 139.175 159.220 139.505 159.690 ;
        RECT 139.675 159.400 139.845 159.860 ;
        RECT 140.015 159.220 140.345 159.690 ;
        RECT 140.515 159.395 140.765 159.860 ;
        RECT 139.175 159.040 140.780 159.220 ;
        RECT 137.335 158.840 137.665 158.870 ;
        RECT 137.110 158.670 137.665 158.840 ;
        RECT 137.335 158.620 137.665 158.670 ;
        RECT 137.835 158.620 140.345 158.870 ;
        RECT 137.835 158.460 138.085 158.620 ;
        RECT 137.355 157.310 137.585 158.450 ;
        RECT 137.755 157.480 138.085 158.460 ;
        RECT 140.515 158.450 140.780 159.040 ;
        RECT 138.255 157.310 138.465 158.450 ;
        RECT 138.740 157.310 139.005 158.450 ;
        RECT 139.175 158.280 140.780 158.450 ;
        RECT 139.175 157.480 139.505 158.280 ;
        RECT 140.015 158.260 140.780 158.280 ;
        RECT 139.675 157.310 139.845 158.110 ;
        RECT 140.015 157.480 140.345 158.260 ;
        RECT 140.515 157.310 140.725 157.770 ;
        RECT 137.230 157.140 140.910 157.310 ;
        RECT 137.415 156.680 137.625 157.140 ;
        RECT 137.795 156.190 138.125 156.970 ;
        RECT 138.295 156.340 138.465 157.140 ;
        RECT 137.360 156.170 138.125 156.190 ;
        RECT 138.635 156.170 138.965 156.970 ;
        RECT 137.360 156.000 138.965 156.170 ;
        RECT 139.135 156.000 139.400 157.140 ;
        RECT 137.360 155.410 137.625 156.000 ;
        RECT 139.880 155.975 140.525 157.140 ;
        RECT 137.795 155.580 139.425 155.830 ;
        RECT 137.360 155.230 138.965 155.410 ;
        RECT 137.375 154.590 137.625 155.055 ;
        RECT 137.795 154.760 138.125 155.230 ;
        RECT 138.295 154.590 138.465 155.050 ;
        RECT 138.635 154.760 138.965 155.230 ;
        RECT 139.135 154.590 139.400 155.050 ;
        RECT 137.230 154.460 139.530 154.590 ;
        RECT 130.390 154.290 136.860 154.460 ;
        RECT 137.225 154.420 139.530 154.460 ;
        RECT 137.225 154.290 139.415 154.420 ;
        RECT 123.640 153.930 130.060 154.100 ;
        RECT 86.690 149.520 118.580 149.690 ;
        RECT 7.290 142.735 35.790 142.915 ;
        RECT 7.290 142.565 35.915 142.735 ;
        RECT 7.290 133.425 7.690 142.565 ;
        RECT 8.265 142.050 8.615 142.220 ;
        RECT 8.905 142.050 9.255 142.220 ;
        RECT 9.545 142.050 9.895 142.220 ;
        RECT 10.185 142.050 10.535 142.220 ;
        RECT 10.825 142.050 11.175 142.220 ;
        RECT 11.465 142.050 11.815 142.220 ;
        RECT 12.105 142.050 12.455 142.220 ;
        RECT 12.745 142.050 13.095 142.220 ;
        RECT 13.385 142.050 13.735 142.220 ;
        RECT 14.025 142.050 14.375 142.220 ;
        RECT 14.665 142.050 15.015 142.220 ;
        RECT 15.305 142.050 15.655 142.220 ;
        RECT 15.945 142.050 16.295 142.220 ;
        RECT 16.585 142.050 16.935 142.220 ;
        RECT 17.225 142.050 17.575 142.220 ;
        RECT 17.865 142.050 18.215 142.220 ;
        RECT 18.505 142.050 18.855 142.220 ;
        RECT 19.145 142.050 19.495 142.220 ;
        RECT 19.785 142.050 20.135 142.220 ;
        RECT 20.425 142.050 20.775 142.220 ;
        RECT 21.065 142.050 21.415 142.220 ;
        RECT 21.705 142.050 22.055 142.220 ;
        RECT 22.345 142.050 22.695 142.220 ;
        RECT 22.985 142.050 23.335 142.220 ;
        RECT 23.625 142.050 23.975 142.220 ;
        RECT 24.265 142.050 24.615 142.220 ;
        RECT 24.905 142.050 25.255 142.220 ;
        RECT 25.545 142.050 25.895 142.220 ;
        RECT 26.185 142.050 26.535 142.220 ;
        RECT 26.825 142.050 27.175 142.220 ;
        RECT 27.465 142.050 27.815 142.220 ;
        RECT 28.690 142.050 29.040 142.220 ;
        RECT 29.900 142.050 30.250 142.220 ;
        RECT 31.110 142.050 31.460 142.220 ;
        RECT 32.320 142.050 32.670 142.220 ;
        RECT 33.530 142.050 33.880 142.220 ;
        RECT 34.740 142.050 35.090 142.220 ;
        RECT 8.035 133.795 8.205 141.835 ;
        RECT 8.675 133.795 8.845 141.835 ;
        RECT 9.315 133.795 9.485 141.835 ;
        RECT 9.955 133.795 10.125 141.835 ;
        RECT 10.595 133.795 10.765 141.835 ;
        RECT 11.235 133.795 11.405 141.835 ;
        RECT 11.875 133.795 12.045 141.835 ;
        RECT 12.515 133.795 12.685 141.835 ;
        RECT 13.155 133.795 13.325 141.835 ;
        RECT 13.795 133.795 13.965 141.835 ;
        RECT 14.435 133.795 14.605 141.835 ;
        RECT 15.075 133.795 15.245 141.835 ;
        RECT 15.715 133.795 15.885 141.835 ;
        RECT 16.355 133.795 16.525 141.835 ;
        RECT 16.995 133.795 17.165 141.835 ;
        RECT 17.635 133.795 17.805 141.835 ;
        RECT 18.275 133.795 18.445 141.835 ;
        RECT 18.915 133.795 19.085 141.835 ;
        RECT 19.555 133.795 19.725 141.835 ;
        RECT 20.195 133.795 20.365 141.835 ;
        RECT 20.835 133.795 21.005 141.835 ;
        RECT 21.475 133.795 21.645 141.835 ;
        RECT 22.115 133.795 22.285 141.835 ;
        RECT 22.755 133.795 22.925 141.835 ;
        RECT 23.395 133.795 23.565 141.835 ;
        RECT 24.035 133.795 24.205 141.835 ;
        RECT 24.675 133.795 24.845 141.835 ;
        RECT 25.315 133.795 25.485 141.835 ;
        RECT 25.955 133.795 26.125 141.835 ;
        RECT 26.595 133.795 26.765 141.835 ;
        RECT 27.235 133.795 27.405 141.835 ;
        RECT 27.875 133.795 28.045 141.835 ;
        RECT 28.460 137.795 28.630 141.835 ;
        RECT 29.100 137.795 29.270 141.835 ;
        RECT 29.670 137.795 29.840 141.835 ;
        RECT 30.310 137.795 30.480 141.835 ;
        RECT 30.880 137.795 31.050 141.835 ;
        RECT 31.520 137.795 31.690 141.835 ;
        RECT 32.090 137.795 32.260 141.835 ;
        RECT 32.730 137.795 32.900 141.835 ;
        RECT 33.300 137.795 33.470 141.835 ;
        RECT 33.940 137.795 34.110 141.835 ;
        RECT 34.510 137.795 34.680 141.835 ;
        RECT 35.150 137.795 35.320 141.835 ;
        RECT 35.745 133.425 35.915 142.565 ;
        RECT 7.290 133.255 35.915 133.425 ;
        RECT 36.090 142.565 75.290 142.915 ;
        RECT 36.090 133.425 36.455 142.565 ;
        RECT 37.495 141.965 37.825 142.135 ;
        RECT 38.455 141.965 38.785 142.135 ;
        RECT 39.415 141.965 39.745 142.135 ;
        RECT 40.375 141.965 40.705 142.135 ;
        RECT 41.335 141.965 41.665 142.135 ;
        RECT 42.295 141.965 42.625 142.135 ;
        RECT 43.255 141.965 43.585 142.135 ;
        RECT 44.125 141.995 44.455 142.165 ;
        RECT 45.260 141.965 45.590 142.135 ;
        RECT 46.130 141.995 46.460 142.165 ;
        RECT 47.340 141.965 47.670 142.135 ;
        RECT 48.300 141.965 48.630 142.135 ;
        RECT 49.260 141.965 49.590 142.135 ;
        RECT 50.220 141.965 50.550 142.135 ;
        RECT 51.180 141.965 51.510 142.135 ;
        RECT 52.140 141.965 52.470 142.135 ;
        RECT 53.100 141.965 53.430 142.135 ;
        RECT 54.060 141.965 54.390 142.135 ;
        RECT 55.020 141.965 55.350 142.135 ;
        RECT 55.980 141.965 56.310 142.135 ;
        RECT 56.940 141.965 57.270 142.135 ;
        RECT 57.900 141.965 58.230 142.135 ;
        RECT 58.940 141.965 59.270 142.135 ;
        RECT 59.900 141.965 60.230 142.135 ;
        RECT 60.460 141.965 60.790 142.135 ;
        RECT 61.510 141.965 61.840 142.135 ;
        RECT 62.555 141.965 62.885 142.135 ;
        RECT 63.610 141.965 63.940 142.135 ;
        RECT 64.655 141.965 64.985 142.135 ;
        RECT 72.950 142.100 73.280 142.270 ;
        RECT 36.855 133.755 37.025 141.795 ;
        RECT 37.335 133.755 37.505 141.795 ;
        RECT 37.815 133.755 37.985 141.795 ;
        RECT 38.295 133.755 38.465 141.795 ;
        RECT 38.775 133.755 38.945 141.795 ;
        RECT 39.255 133.755 39.425 141.795 ;
        RECT 39.735 133.755 39.905 141.795 ;
        RECT 40.215 133.755 40.385 141.795 ;
        RECT 40.695 133.755 40.865 141.795 ;
        RECT 41.175 133.755 41.345 141.795 ;
        RECT 41.655 133.755 41.825 141.795 ;
        RECT 42.135 133.755 42.305 141.795 ;
        RECT 42.615 133.755 42.785 141.795 ;
        RECT 43.095 133.755 43.265 141.795 ;
        RECT 43.575 133.755 43.745 141.795 ;
        RECT 44.055 133.755 44.225 141.795 ;
        RECT 44.620 133.755 44.790 141.795 ;
        RECT 45.100 133.755 45.270 141.795 ;
        RECT 45.580 133.755 45.750 141.795 ;
        RECT 46.060 133.755 46.230 141.795 ;
        RECT 46.700 133.755 46.870 141.795 ;
        RECT 47.180 133.755 47.350 141.795 ;
        RECT 47.660 133.755 47.830 141.795 ;
        RECT 48.140 133.755 48.310 141.795 ;
        RECT 48.620 133.755 48.790 141.795 ;
        RECT 49.100 133.755 49.270 141.795 ;
        RECT 49.580 133.755 49.750 141.795 ;
        RECT 50.060 133.755 50.230 141.795 ;
        RECT 50.540 133.755 50.710 141.795 ;
        RECT 51.020 133.755 51.190 141.795 ;
        RECT 51.500 133.755 51.670 141.795 ;
        RECT 51.980 133.755 52.150 141.795 ;
        RECT 52.460 133.755 52.630 141.795 ;
        RECT 52.940 133.755 53.110 141.795 ;
        RECT 53.420 133.755 53.590 141.795 ;
        RECT 53.900 133.755 54.070 141.795 ;
        RECT 54.380 133.755 54.550 141.795 ;
        RECT 54.860 133.755 55.030 141.795 ;
        RECT 55.340 133.755 55.510 141.795 ;
        RECT 55.820 133.755 55.990 141.795 ;
        RECT 56.300 133.755 56.470 141.795 ;
        RECT 56.780 133.755 56.950 141.795 ;
        RECT 57.260 133.755 57.430 141.795 ;
        RECT 57.740 133.755 57.910 141.795 ;
        RECT 58.300 139.755 58.470 141.795 ;
        RECT 58.780 139.755 58.950 141.795 ;
        RECT 59.260 139.755 59.430 141.795 ;
        RECT 59.740 139.755 59.910 141.795 ;
        RECT 60.300 139.755 60.470 141.795 ;
        RECT 60.780 139.755 60.950 141.795 ;
        RECT 61.350 139.755 61.520 141.795 ;
        RECT 61.830 139.755 62.000 141.795 ;
        RECT 62.400 139.755 62.570 141.795 ;
        RECT 62.880 139.755 63.050 141.795 ;
        RECT 63.450 139.755 63.620 141.795 ;
        RECT 63.930 139.755 64.100 141.795 ;
        RECT 64.500 139.755 64.670 141.795 ;
        RECT 64.980 139.755 65.150 141.795 ;
        RECT 72.790 140.890 72.960 141.930 ;
        RECT 73.270 140.890 73.440 141.930 ;
        RECT 72.950 140.085 73.280 140.255 ;
        RECT 72.790 138.875 72.960 139.915 ;
        RECT 73.270 138.875 73.440 139.915 ;
        RECT 72.960 137.920 73.290 138.090 ;
        RECT 72.800 136.710 72.970 137.750 ;
        RECT 73.280 136.710 73.450 137.750 ;
        RECT 58.940 135.965 59.270 136.135 ;
        RECT 59.900 135.965 60.230 136.135 ;
        RECT 60.455 135.965 60.785 136.135 ;
        RECT 61.510 135.965 61.840 136.135 ;
        RECT 62.560 135.965 62.890 136.135 ;
        RECT 63.610 135.965 63.940 136.135 ;
        RECT 64.655 135.985 64.985 136.155 ;
        RECT 65.710 135.965 66.040 136.135 ;
        RECT 67.240 135.970 67.570 136.140 ;
        RECT 68.200 135.970 68.530 136.140 ;
        RECT 68.760 135.970 69.090 136.140 ;
        RECT 69.810 135.970 70.140 136.140 ;
        RECT 70.860 135.970 71.190 136.140 ;
        RECT 71.910 135.970 72.240 136.140 ;
        RECT 72.960 135.970 73.290 136.140 ;
        RECT 58.300 133.755 58.470 135.795 ;
        RECT 58.780 133.755 58.950 135.795 ;
        RECT 59.260 133.755 59.430 135.795 ;
        RECT 59.740 133.755 59.910 135.795 ;
        RECT 60.300 133.755 60.470 135.795 ;
        RECT 60.780 133.755 60.950 135.795 ;
        RECT 61.350 133.755 61.520 135.795 ;
        RECT 61.830 133.755 62.000 135.795 ;
        RECT 62.400 133.755 62.570 135.795 ;
        RECT 62.880 133.755 63.050 135.795 ;
        RECT 63.450 133.755 63.620 135.795 ;
        RECT 63.930 133.755 64.100 135.795 ;
        RECT 64.500 133.755 64.670 135.795 ;
        RECT 64.980 133.755 65.150 135.795 ;
        RECT 65.550 133.755 65.720 135.795 ;
        RECT 66.030 133.755 66.200 135.795 ;
        RECT 66.600 133.760 66.770 135.800 ;
        RECT 67.080 133.760 67.250 135.800 ;
        RECT 67.560 133.760 67.730 135.800 ;
        RECT 68.040 133.760 68.210 135.800 ;
        RECT 68.600 134.760 68.770 135.800 ;
        RECT 69.080 134.760 69.250 135.800 ;
        RECT 69.650 134.760 69.820 135.800 ;
        RECT 70.130 134.760 70.300 135.800 ;
        RECT 70.700 134.760 70.870 135.800 ;
        RECT 71.180 134.760 71.350 135.800 ;
        RECT 71.750 134.760 71.920 135.800 ;
        RECT 72.230 134.760 72.400 135.800 ;
        RECT 72.800 134.760 72.970 135.800 ;
        RECT 73.280 134.760 73.450 135.800 ;
        RECT 74.975 133.425 75.290 142.565 ;
        RECT 7.290 133.065 35.590 133.255 ;
        RECT 36.090 133.065 75.290 133.425 ;
        RECT 85.825 142.565 125.025 142.915 ;
        RECT 125.325 142.735 153.825 142.915 ;
        RECT 85.825 133.425 86.140 142.565 ;
        RECT 87.835 142.100 88.165 142.270 ;
        RECT 96.130 141.965 96.460 142.135 ;
        RECT 97.175 141.965 97.505 142.135 ;
        RECT 98.230 141.965 98.560 142.135 ;
        RECT 99.275 141.965 99.605 142.135 ;
        RECT 100.325 141.965 100.655 142.135 ;
        RECT 100.885 141.965 101.215 142.135 ;
        RECT 101.845 141.965 102.175 142.135 ;
        RECT 102.885 141.965 103.215 142.135 ;
        RECT 103.845 141.965 104.175 142.135 ;
        RECT 104.805 141.965 105.135 142.135 ;
        RECT 105.765 141.965 106.095 142.135 ;
        RECT 106.725 141.965 107.055 142.135 ;
        RECT 107.685 141.965 108.015 142.135 ;
        RECT 108.645 141.965 108.975 142.135 ;
        RECT 109.605 141.965 109.935 142.135 ;
        RECT 110.565 141.965 110.895 142.135 ;
        RECT 111.525 141.965 111.855 142.135 ;
        RECT 112.485 141.965 112.815 142.135 ;
        RECT 113.445 141.965 113.775 142.135 ;
        RECT 114.655 141.995 114.985 142.165 ;
        RECT 115.525 141.965 115.855 142.135 ;
        RECT 116.660 141.995 116.990 142.165 ;
        RECT 117.530 141.965 117.860 142.135 ;
        RECT 118.490 141.965 118.820 142.135 ;
        RECT 119.450 141.965 119.780 142.135 ;
        RECT 120.410 141.965 120.740 142.135 ;
        RECT 121.370 141.965 121.700 142.135 ;
        RECT 122.330 141.965 122.660 142.135 ;
        RECT 123.290 141.965 123.620 142.135 ;
        RECT 87.675 140.890 87.845 141.930 ;
        RECT 88.155 140.890 88.325 141.930 ;
        RECT 87.835 140.085 88.165 140.255 ;
        RECT 87.675 138.875 87.845 139.915 ;
        RECT 88.155 138.875 88.325 139.915 ;
        RECT 95.965 139.755 96.135 141.795 ;
        RECT 96.445 139.755 96.615 141.795 ;
        RECT 97.015 139.755 97.185 141.795 ;
        RECT 97.495 139.755 97.665 141.795 ;
        RECT 98.065 139.755 98.235 141.795 ;
        RECT 98.545 139.755 98.715 141.795 ;
        RECT 99.115 139.755 99.285 141.795 ;
        RECT 99.595 139.755 99.765 141.795 ;
        RECT 100.165 139.755 100.335 141.795 ;
        RECT 100.645 139.755 100.815 141.795 ;
        RECT 101.205 139.755 101.375 141.795 ;
        RECT 101.685 139.755 101.855 141.795 ;
        RECT 102.165 139.755 102.335 141.795 ;
        RECT 102.645 139.755 102.815 141.795 ;
        RECT 87.825 137.920 88.155 138.090 ;
        RECT 87.665 136.710 87.835 137.750 ;
        RECT 88.145 136.710 88.315 137.750 ;
        RECT 87.825 135.970 88.155 136.140 ;
        RECT 88.875 135.970 89.205 136.140 ;
        RECT 89.925 135.970 90.255 136.140 ;
        RECT 90.975 135.970 91.305 136.140 ;
        RECT 92.025 135.970 92.355 136.140 ;
        RECT 92.585 135.970 92.915 136.140 ;
        RECT 93.545 135.970 93.875 136.140 ;
        RECT 95.075 135.965 95.405 136.135 ;
        RECT 96.130 135.985 96.460 136.155 ;
        RECT 97.175 135.965 97.505 136.135 ;
        RECT 98.225 135.965 98.555 136.135 ;
        RECT 99.275 135.965 99.605 136.135 ;
        RECT 100.330 135.965 100.660 136.135 ;
        RECT 100.885 135.965 101.215 136.135 ;
        RECT 101.845 135.965 102.175 136.135 ;
        RECT 87.665 134.760 87.835 135.800 ;
        RECT 88.145 134.760 88.315 135.800 ;
        RECT 88.715 134.760 88.885 135.800 ;
        RECT 89.195 134.760 89.365 135.800 ;
        RECT 89.765 134.760 89.935 135.800 ;
        RECT 90.245 134.760 90.415 135.800 ;
        RECT 90.815 134.760 90.985 135.800 ;
        RECT 91.295 134.760 91.465 135.800 ;
        RECT 91.865 134.760 92.035 135.800 ;
        RECT 92.345 134.760 92.515 135.800 ;
        RECT 92.905 133.760 93.075 135.800 ;
        RECT 93.385 133.760 93.555 135.800 ;
        RECT 93.865 133.760 94.035 135.800 ;
        RECT 94.345 133.760 94.515 135.800 ;
        RECT 94.915 133.755 95.085 135.795 ;
        RECT 95.395 133.755 95.565 135.795 ;
        RECT 95.965 133.755 96.135 135.795 ;
        RECT 96.445 133.755 96.615 135.795 ;
        RECT 97.015 133.755 97.185 135.795 ;
        RECT 97.495 133.755 97.665 135.795 ;
        RECT 98.065 133.755 98.235 135.795 ;
        RECT 98.545 133.755 98.715 135.795 ;
        RECT 99.115 133.755 99.285 135.795 ;
        RECT 99.595 133.755 99.765 135.795 ;
        RECT 100.165 133.755 100.335 135.795 ;
        RECT 100.645 133.755 100.815 135.795 ;
        RECT 101.205 133.755 101.375 135.795 ;
        RECT 101.685 133.755 101.855 135.795 ;
        RECT 102.165 133.755 102.335 135.795 ;
        RECT 102.645 133.755 102.815 135.795 ;
        RECT 103.205 133.755 103.375 141.795 ;
        RECT 103.685 133.755 103.855 141.795 ;
        RECT 104.165 133.755 104.335 141.795 ;
        RECT 104.645 133.755 104.815 141.795 ;
        RECT 105.125 133.755 105.295 141.795 ;
        RECT 105.605 133.755 105.775 141.795 ;
        RECT 106.085 133.755 106.255 141.795 ;
        RECT 106.565 133.755 106.735 141.795 ;
        RECT 107.045 133.755 107.215 141.795 ;
        RECT 107.525 133.755 107.695 141.795 ;
        RECT 108.005 133.755 108.175 141.795 ;
        RECT 108.485 133.755 108.655 141.795 ;
        RECT 108.965 133.755 109.135 141.795 ;
        RECT 109.445 133.755 109.615 141.795 ;
        RECT 109.925 133.755 110.095 141.795 ;
        RECT 110.405 133.755 110.575 141.795 ;
        RECT 110.885 133.755 111.055 141.795 ;
        RECT 111.365 133.755 111.535 141.795 ;
        RECT 111.845 133.755 112.015 141.795 ;
        RECT 112.325 133.755 112.495 141.795 ;
        RECT 112.805 133.755 112.975 141.795 ;
        RECT 113.285 133.755 113.455 141.795 ;
        RECT 113.765 133.755 113.935 141.795 ;
        RECT 114.245 133.755 114.415 141.795 ;
        RECT 114.885 133.755 115.055 141.795 ;
        RECT 115.365 133.755 115.535 141.795 ;
        RECT 115.845 133.755 116.015 141.795 ;
        RECT 116.325 133.755 116.495 141.795 ;
        RECT 116.890 133.755 117.060 141.795 ;
        RECT 117.370 133.755 117.540 141.795 ;
        RECT 117.850 133.755 118.020 141.795 ;
        RECT 118.330 133.755 118.500 141.795 ;
        RECT 118.810 133.755 118.980 141.795 ;
        RECT 119.290 133.755 119.460 141.795 ;
        RECT 119.770 133.755 119.940 141.795 ;
        RECT 120.250 133.755 120.420 141.795 ;
        RECT 120.730 133.755 120.900 141.795 ;
        RECT 121.210 133.755 121.380 141.795 ;
        RECT 121.690 133.755 121.860 141.795 ;
        RECT 122.170 133.755 122.340 141.795 ;
        RECT 122.650 133.755 122.820 141.795 ;
        RECT 123.130 133.755 123.300 141.795 ;
        RECT 123.610 133.755 123.780 141.795 ;
        RECT 124.090 133.755 124.260 141.795 ;
        RECT 124.660 133.425 125.025 142.565 ;
        RECT 85.825 133.065 125.025 133.425 ;
        RECT 125.200 142.565 153.825 142.735 ;
        RECT 125.200 133.425 125.370 142.565 ;
        RECT 126.025 142.050 126.375 142.220 ;
        RECT 127.235 142.050 127.585 142.220 ;
        RECT 128.445 142.050 128.795 142.220 ;
        RECT 129.655 142.050 130.005 142.220 ;
        RECT 130.865 142.050 131.215 142.220 ;
        RECT 132.075 142.050 132.425 142.220 ;
        RECT 133.300 142.050 133.650 142.220 ;
        RECT 133.940 142.050 134.290 142.220 ;
        RECT 134.580 142.050 134.930 142.220 ;
        RECT 135.220 142.050 135.570 142.220 ;
        RECT 135.860 142.050 136.210 142.220 ;
        RECT 136.500 142.050 136.850 142.220 ;
        RECT 137.140 142.050 137.490 142.220 ;
        RECT 137.780 142.050 138.130 142.220 ;
        RECT 138.420 142.050 138.770 142.220 ;
        RECT 139.060 142.050 139.410 142.220 ;
        RECT 139.700 142.050 140.050 142.220 ;
        RECT 140.340 142.050 140.690 142.220 ;
        RECT 140.980 142.050 141.330 142.220 ;
        RECT 141.620 142.050 141.970 142.220 ;
        RECT 142.260 142.050 142.610 142.220 ;
        RECT 142.900 142.050 143.250 142.220 ;
        RECT 143.540 142.050 143.890 142.220 ;
        RECT 144.180 142.050 144.530 142.220 ;
        RECT 144.820 142.050 145.170 142.220 ;
        RECT 145.460 142.050 145.810 142.220 ;
        RECT 146.100 142.050 146.450 142.220 ;
        RECT 146.740 142.050 147.090 142.220 ;
        RECT 147.380 142.050 147.730 142.220 ;
        RECT 148.020 142.050 148.370 142.220 ;
        RECT 148.660 142.050 149.010 142.220 ;
        RECT 149.300 142.050 149.650 142.220 ;
        RECT 149.940 142.050 150.290 142.220 ;
        RECT 150.580 142.050 150.930 142.220 ;
        RECT 151.220 142.050 151.570 142.220 ;
        RECT 151.860 142.050 152.210 142.220 ;
        RECT 152.500 142.050 152.850 142.220 ;
        RECT 125.795 137.795 125.965 141.835 ;
        RECT 126.435 137.795 126.605 141.835 ;
        RECT 127.005 137.795 127.175 141.835 ;
        RECT 127.645 137.795 127.815 141.835 ;
        RECT 128.215 137.795 128.385 141.835 ;
        RECT 128.855 137.795 129.025 141.835 ;
        RECT 129.425 137.795 129.595 141.835 ;
        RECT 130.065 137.795 130.235 141.835 ;
        RECT 130.635 137.795 130.805 141.835 ;
        RECT 131.275 137.795 131.445 141.835 ;
        RECT 131.845 137.795 132.015 141.835 ;
        RECT 132.485 137.795 132.655 141.835 ;
        RECT 133.070 133.795 133.240 141.835 ;
        RECT 133.710 133.795 133.880 141.835 ;
        RECT 134.350 133.795 134.520 141.835 ;
        RECT 134.990 133.795 135.160 141.835 ;
        RECT 135.630 133.795 135.800 141.835 ;
        RECT 136.270 133.795 136.440 141.835 ;
        RECT 136.910 133.795 137.080 141.835 ;
        RECT 137.550 133.795 137.720 141.835 ;
        RECT 138.190 133.795 138.360 141.835 ;
        RECT 138.830 133.795 139.000 141.835 ;
        RECT 139.470 133.795 139.640 141.835 ;
        RECT 140.110 133.795 140.280 141.835 ;
        RECT 140.750 133.795 140.920 141.835 ;
        RECT 141.390 133.795 141.560 141.835 ;
        RECT 142.030 133.795 142.200 141.835 ;
        RECT 142.670 133.795 142.840 141.835 ;
        RECT 143.310 133.795 143.480 141.835 ;
        RECT 143.950 133.795 144.120 141.835 ;
        RECT 144.590 133.795 144.760 141.835 ;
        RECT 145.230 133.795 145.400 141.835 ;
        RECT 145.870 133.795 146.040 141.835 ;
        RECT 146.510 133.795 146.680 141.835 ;
        RECT 147.150 133.795 147.320 141.835 ;
        RECT 147.790 133.795 147.960 141.835 ;
        RECT 148.430 133.795 148.600 141.835 ;
        RECT 149.070 133.795 149.240 141.835 ;
        RECT 149.710 133.795 149.880 141.835 ;
        RECT 150.350 133.795 150.520 141.835 ;
        RECT 150.990 133.795 151.160 141.835 ;
        RECT 151.630 133.795 151.800 141.835 ;
        RECT 152.270 133.795 152.440 141.835 ;
        RECT 152.910 133.795 153.080 141.835 ;
        RECT 153.425 133.425 153.825 142.565 ;
        RECT 125.200 133.255 153.825 133.425 ;
        RECT 125.525 133.065 153.825 133.255 ;
        RECT 7.490 127.290 8.190 127.490 ;
        RECT 152.925 127.290 153.625 127.490 ;
        RECT 7.740 126.040 7.940 127.290 ;
        RECT 73.490 127.040 74.190 127.240 ;
        RECT 86.925 127.040 87.625 127.240 ;
        RECT 73.740 126.040 73.940 127.040 ;
        RECT 6.990 5.940 7.190 126.040 ;
        RECT 7.360 125.940 73.940 126.040 ;
        RECT 87.175 126.040 87.375 127.040 ;
        RECT 153.175 126.040 153.375 127.290 ;
        RECT 87.175 125.940 153.755 126.040 ;
        RECT 7.360 125.840 73.920 125.940 ;
        RECT 87.195 125.840 153.755 125.940 ;
        RECT 153.925 5.940 154.125 126.040 ;
        RECT 7.360 5.590 73.920 5.790 ;
        RECT 87.195 5.590 153.755 5.790 ;
      LAYER met1 ;
        RECT 98.540 220.080 98.940 220.140 ;
        RECT 98.540 219.940 150.210 220.080 ;
        RECT 98.540 219.840 98.940 219.940 ;
        RECT 99.490 219.735 99.810 219.795 ;
        RECT 143.190 219.735 143.510 219.795 ;
        RECT 10.215 219.240 10.515 219.640 ;
        RECT 99.490 219.595 143.510 219.735 ;
        RECT 99.490 219.535 99.810 219.595 ;
        RECT 143.190 219.535 143.510 219.595 ;
        RECT 9.815 217.940 10.115 218.340 ;
        RECT 9.465 216.590 9.765 216.990 ;
        RECT 9.165 215.190 9.465 215.590 ;
        RECT 8.865 213.840 9.165 214.240 ;
        RECT 8.565 212.440 8.865 212.840 ;
        RECT 8.265 211.140 8.565 211.540 ;
        RECT 7.965 209.790 8.265 210.190 ;
        RECT 7.665 208.390 7.965 208.790 ;
        RECT 7.365 207.040 7.665 207.440 ;
        RECT 7.065 205.740 7.365 206.140 ;
        RECT 6.765 204.340 7.065 204.740 ;
        RECT 6.465 202.990 6.765 203.390 ;
        RECT 6.165 201.590 6.465 201.990 ;
        RECT 5.865 200.290 6.165 200.690 ;
        RECT 5.565 198.940 5.865 199.340 ;
        RECT 5.265 197.590 5.565 197.990 ;
        RECT 4.965 196.140 5.265 196.540 ;
        RECT 4.665 194.790 4.965 195.190 ;
        RECT 4.365 193.490 4.665 193.890 ;
        RECT 4.065 192.040 4.365 192.440 ;
        RECT 3.765 190.690 4.065 191.090 ;
        RECT 3.465 189.290 3.765 189.690 ;
        RECT 3.615 168.075 3.765 189.290 ;
        RECT 3.915 180.015 4.065 190.690 ;
        RECT 4.215 180.315 4.365 192.040 ;
        RECT 4.515 180.615 4.665 193.490 ;
        RECT 4.815 180.915 4.965 194.790 ;
        RECT 5.115 181.215 5.265 196.140 ;
        RECT 5.415 181.515 5.565 197.590 ;
        RECT 5.715 181.810 5.865 198.940 ;
        RECT 6.015 182.115 6.165 200.290 ;
        RECT 6.315 182.415 6.465 201.590 ;
        RECT 6.615 182.715 6.765 202.990 ;
        RECT 6.915 183.140 7.065 204.340 ;
        RECT 7.215 183.440 7.365 205.740 ;
        RECT 7.515 183.740 7.665 207.040 ;
        RECT 7.815 184.040 7.965 208.390 ;
        RECT 8.115 184.340 8.265 209.790 ;
        RECT 8.415 184.640 8.565 211.140 ;
        RECT 8.715 184.940 8.865 212.440 ;
        RECT 9.015 185.240 9.165 213.840 ;
        RECT 9.315 185.540 9.465 215.190 ;
        RECT 9.615 185.840 9.765 216.590 ;
        RECT 9.915 186.140 10.065 217.940 ;
        RECT 10.365 186.465 10.515 219.240 ;
        RECT 45.670 219.395 45.990 219.455 ;
        RECT 145.030 219.395 145.350 219.455 ;
        RECT 45.670 219.255 145.350 219.395 ;
        RECT 45.670 219.195 45.990 219.255 ;
        RECT 145.030 219.195 145.350 219.255 ;
        RECT 59.930 219.055 60.250 219.115 ;
        RECT 133.530 219.055 133.850 219.115 ;
        RECT 59.930 218.915 133.850 219.055 ;
        RECT 59.930 218.855 60.250 218.915 ;
        RECT 133.530 218.855 133.850 218.915 ;
        RECT 43.370 218.715 43.690 218.775 ;
        RECT 49.350 218.715 49.670 218.775 ;
        RECT 64.990 218.715 65.310 218.775 ;
        RECT 43.370 218.575 65.310 218.715 ;
        RECT 43.370 218.515 43.690 218.575 ;
        RECT 49.350 218.515 49.670 218.575 ;
        RECT 64.990 218.515 65.310 218.575 ;
        RECT 84.310 218.715 84.630 218.775 ;
        RECT 110.530 218.715 110.850 218.775 ;
        RECT 84.310 218.575 110.850 218.715 ;
        RECT 84.310 218.515 84.630 218.575 ;
        RECT 110.530 218.515 110.850 218.575 ;
        RECT 14.390 218.375 14.710 218.435 ;
        RECT 21.750 218.375 22.070 218.435 ;
        RECT 14.390 218.235 22.070 218.375 ;
        RECT 14.390 218.175 14.710 218.235 ;
        RECT 21.750 218.175 22.070 218.235 ;
        RECT 22.670 218.375 22.990 218.435 ;
        RECT 98.110 218.375 98.430 218.435 ;
        RECT 22.670 218.235 98.430 218.375 ;
        RECT 22.670 218.175 22.990 218.235 ;
        RECT 98.110 218.175 98.430 218.235 ;
        RECT 103.170 218.375 103.490 218.435 ;
        RECT 140.890 218.375 141.210 218.435 ;
        RECT 103.170 218.235 141.210 218.375 ;
        RECT 103.170 218.175 103.490 218.235 ;
        RECT 140.890 218.175 141.210 218.235 ;
        RECT 13.860 217.555 147.720 218.035 ;
        RECT 13.930 217.355 14.250 217.415 ;
        RECT 18.545 217.355 18.835 217.400 ;
        RECT 13.930 217.215 18.835 217.355 ;
        RECT 13.930 217.155 14.250 217.215 ;
        RECT 18.545 217.170 18.835 217.215 ;
        RECT 22.670 217.155 22.990 217.415 ;
        RECT 27.285 217.170 27.575 217.400 ;
        RECT 29.125 217.355 29.415 217.400 ;
        RECT 29.125 217.215 38.540 217.355 ;
        RECT 29.125 217.170 29.415 217.215 ;
        RECT 14.850 217.015 15.170 217.075 ;
        RECT 15.325 217.015 15.615 217.060 ;
        RECT 14.850 216.875 15.615 217.015 ;
        RECT 14.850 216.815 15.170 216.875 ;
        RECT 15.325 216.830 15.615 216.875 ;
        RECT 17.165 217.015 17.455 217.060 ;
        RECT 22.210 217.015 22.530 217.075 ;
        RECT 17.165 216.875 22.530 217.015 ;
        RECT 17.165 216.830 17.455 216.875 ;
        RECT 22.210 216.815 22.530 216.875 ;
        RECT 19.465 216.490 19.755 216.720 ;
        RECT 19.540 216.335 19.680 216.490 ;
        RECT 21.290 216.475 21.610 216.735 ;
        RECT 21.750 216.475 22.070 216.735 ;
        RECT 26.365 216.675 26.655 216.720 ;
        RECT 27.360 216.675 27.500 217.170 ;
        RECT 36.025 217.015 36.315 217.060 ;
        RECT 37.405 217.015 37.695 217.060 ;
        RECT 26.365 216.535 27.500 216.675 ;
        RECT 29.200 216.875 35.780 217.015 ;
        RECT 26.365 216.490 26.655 216.535 ;
        RECT 29.200 216.335 29.340 216.875 ;
        RECT 29.585 216.675 29.875 216.720 ;
        RECT 31.410 216.675 31.730 216.735 ;
        RECT 29.585 216.535 31.730 216.675 ;
        RECT 29.585 216.490 29.875 216.535 ;
        RECT 31.410 216.475 31.730 216.535 ;
        RECT 31.870 216.475 32.190 216.735 ;
        RECT 19.540 216.195 29.340 216.335 ;
        RECT 30.030 216.335 30.350 216.395 ;
        RECT 30.505 216.335 30.795 216.380 ;
        RECT 30.030 216.195 35.320 216.335 ;
        RECT 30.030 216.135 30.350 216.195 ;
        RECT 30.505 216.150 30.795 216.195 ;
        RECT 25.905 215.995 26.195 216.040 ;
        RECT 31.870 215.995 32.190 216.055 ;
        RECT 25.905 215.855 32.190 215.995 ;
        RECT 25.905 215.810 26.195 215.855 ;
        RECT 31.870 215.795 32.190 215.855 ;
        RECT 20.370 215.455 20.690 215.715 ;
        RECT 26.810 215.655 27.130 215.715 ;
        RECT 32.345 215.655 32.635 215.700 ;
        RECT 26.810 215.515 32.635 215.655 ;
        RECT 35.180 215.655 35.320 216.195 ;
        RECT 35.640 215.995 35.780 216.875 ;
        RECT 36.025 216.875 37.695 217.015 ;
        RECT 38.400 217.015 38.540 217.215 ;
        RECT 38.770 217.155 39.090 217.415 ;
        RECT 40.165 217.170 40.455 217.400 ;
        RECT 39.230 217.015 39.550 217.075 ;
        RECT 38.400 216.875 39.550 217.015 ;
        RECT 36.025 216.830 36.315 216.875 ;
        RECT 37.405 216.830 37.695 216.875 ;
        RECT 39.230 216.815 39.550 216.875 ;
        RECT 36.485 216.675 36.775 216.720 ;
        RECT 40.240 216.675 40.380 217.170 ;
        RECT 50.730 217.155 51.050 217.415 ;
        RECT 53.045 217.170 53.335 217.400 ;
        RECT 62.690 217.355 63.010 217.415 ;
        RECT 66.845 217.355 67.135 217.400 ;
        RECT 62.690 217.215 67.135 217.355 ;
        RECT 46.130 216.815 46.450 217.075 ;
        RECT 48.905 217.015 49.195 217.060 ;
        RECT 50.285 217.015 50.575 217.060 ;
        RECT 48.905 216.875 50.575 217.015 ;
        RECT 48.905 216.830 49.195 216.875 ;
        RECT 50.285 216.830 50.575 216.875 ;
        RECT 36.485 216.535 40.380 216.675 ;
        RECT 41.530 216.675 41.850 216.735 ;
        RECT 42.005 216.675 42.295 216.720 ;
        RECT 41.530 216.535 42.295 216.675 ;
        RECT 36.485 216.490 36.775 216.535 ;
        RECT 41.530 216.475 41.850 216.535 ;
        RECT 42.005 216.490 42.295 216.535 ;
        RECT 49.365 216.675 49.655 216.720 ;
        RECT 53.120 216.675 53.260 217.170 ;
        RECT 62.690 217.155 63.010 217.215 ;
        RECT 66.845 217.170 67.135 217.215 ;
        RECT 74.650 217.355 74.970 217.415 ;
        RECT 76.045 217.355 76.335 217.400 ;
        RECT 74.650 217.215 76.335 217.355 ;
        RECT 74.650 217.155 74.970 217.215 ;
        RECT 76.045 217.170 76.335 217.215 ;
        RECT 84.770 217.355 85.090 217.415 ;
        RECT 105.470 217.355 105.790 217.415 ;
        RECT 84.770 217.215 96.040 217.355 ;
        RECT 84.770 217.155 85.090 217.215 ;
        RECT 53.490 217.015 53.810 217.075 ;
        RECT 55.345 217.015 55.635 217.060 ;
        RECT 64.530 217.015 64.850 217.075 ;
        RECT 53.490 216.875 55.635 217.015 ;
        RECT 53.490 216.815 53.810 216.875 ;
        RECT 55.345 216.830 55.635 216.875 ;
        RECT 63.240 216.875 64.850 217.015 ;
        RECT 49.365 216.535 53.260 216.675 ;
        RECT 49.365 216.490 49.655 216.535 ;
        RECT 54.885 216.490 55.175 216.720 ;
        RECT 60.405 216.675 60.695 216.720 ;
        RECT 62.690 216.675 63.010 216.735 ;
        RECT 63.240 216.720 63.380 216.875 ;
        RECT 64.530 216.815 64.850 216.875 ;
        RECT 70.510 217.015 70.830 217.075 ;
        RECT 75.585 217.015 75.875 217.060 ;
        RECT 70.510 216.875 75.875 217.015 ;
        RECT 70.510 216.815 70.830 216.875 ;
        RECT 75.585 216.830 75.875 216.875 ;
        RECT 77.410 217.015 77.730 217.075 ;
        RECT 87.545 217.015 87.835 217.060 ;
        RECT 77.410 216.875 87.835 217.015 ;
        RECT 77.410 216.815 77.730 216.875 ;
        RECT 87.545 216.830 87.835 216.875 ;
        RECT 60.405 216.535 63.010 216.675 ;
        RECT 60.405 216.490 60.695 216.535 ;
        RECT 39.690 216.335 40.010 216.395 ;
        RECT 42.465 216.335 42.755 216.380 ;
        RECT 39.690 216.195 42.755 216.335 ;
        RECT 39.690 216.135 40.010 216.195 ;
        RECT 42.465 216.150 42.755 216.195 ;
        RECT 43.370 216.135 43.690 216.395 ;
        RECT 46.590 216.135 46.910 216.395 ;
        RECT 47.050 216.135 47.370 216.395 ;
        RECT 54.960 215.995 55.100 216.490 ;
        RECT 62.690 216.475 63.010 216.535 ;
        RECT 63.165 216.490 63.455 216.720 ;
        RECT 63.625 216.490 63.915 216.720 ;
        RECT 64.085 216.675 64.375 216.720 ;
        RECT 66.385 216.675 66.675 216.720 ;
        RECT 64.085 216.535 66.675 216.675 ;
        RECT 64.085 216.490 64.375 216.535 ;
        RECT 66.385 216.490 66.675 216.535 ;
        RECT 70.050 216.675 70.370 216.735 ;
        RECT 95.900 216.720 96.040 217.215 ;
        RECT 105.470 217.215 119.500 217.355 ;
        RECT 105.470 217.155 105.790 217.215 ;
        RECT 103.630 217.015 103.950 217.075 ;
        RECT 97.740 216.875 103.950 217.015 ;
        RECT 79.725 216.675 80.015 216.720 ;
        RECT 85.705 216.675 85.995 216.720 ;
        RECT 70.050 216.535 85.995 216.675 ;
        RECT 56.265 216.335 56.555 216.380 ;
        RECT 57.170 216.335 57.490 216.395 ;
        RECT 56.265 216.195 57.490 216.335 ;
        RECT 56.265 216.150 56.555 216.195 ;
        RECT 57.170 216.135 57.490 216.195 ;
        RECT 62.230 216.335 62.550 216.395 ;
        RECT 63.700 216.335 63.840 216.490 ;
        RECT 70.050 216.475 70.370 216.535 ;
        RECT 79.725 216.490 80.015 216.535 ;
        RECT 85.705 216.490 85.995 216.535 ;
        RECT 95.825 216.675 96.115 216.720 ;
        RECT 97.190 216.675 97.510 216.735 ;
        RECT 95.825 216.535 97.510 216.675 ;
        RECT 95.825 216.490 96.115 216.535 ;
        RECT 62.230 216.195 63.840 216.335 ;
        RECT 62.230 216.135 62.550 216.195 ;
        RECT 69.130 216.135 69.450 216.395 ;
        RECT 78.790 216.135 79.110 216.395 ;
        RECT 79.250 216.335 79.570 216.395 ;
        RECT 80.645 216.335 80.935 216.380 ;
        RECT 79.250 216.195 80.935 216.335 ;
        RECT 79.250 216.135 79.570 216.195 ;
        RECT 80.645 216.150 80.935 216.195 ;
        RECT 84.770 216.135 85.090 216.395 ;
        RECT 85.780 216.335 85.920 216.490 ;
        RECT 97.190 216.475 97.510 216.535 ;
        RECT 97.740 216.335 97.880 216.875 ;
        RECT 103.630 216.815 103.950 216.875 ;
        RECT 110.985 217.015 111.635 217.060 ;
        RECT 114.585 217.015 114.875 217.060 ;
        RECT 110.985 216.875 114.875 217.015 ;
        RECT 110.985 216.830 111.635 216.875 ;
        RECT 114.285 216.830 114.875 216.875 ;
        RECT 98.570 216.675 98.890 216.735 ;
        RECT 101.345 216.675 101.635 216.720 ;
        RECT 98.570 216.535 101.635 216.675 ;
        RECT 98.570 216.475 98.890 216.535 ;
        RECT 101.345 216.490 101.635 216.535 ;
        RECT 104.565 216.490 104.855 216.720 ;
        RECT 107.790 216.675 108.080 216.720 ;
        RECT 109.625 216.675 109.915 216.720 ;
        RECT 113.205 216.675 113.495 216.720 ;
        RECT 107.790 216.535 113.495 216.675 ;
        RECT 107.790 216.490 108.080 216.535 ;
        RECT 109.625 216.490 109.915 216.535 ;
        RECT 113.205 216.490 113.495 216.535 ;
        RECT 114.285 216.515 114.575 216.830 ;
        RECT 119.360 216.720 119.500 217.215 ;
        RECT 122.120 217.215 125.480 217.355 ;
        RECT 122.120 216.720 122.260 217.215 ;
        RECT 85.780 216.195 97.880 216.335 ;
        RECT 99.030 216.335 99.350 216.395 ;
        RECT 102.710 216.335 103.030 216.395 ;
        RECT 99.030 216.195 103.030 216.335 ;
        RECT 99.030 216.135 99.350 216.195 ;
        RECT 102.710 216.135 103.030 216.195 ;
        RECT 79.710 215.995 80.030 216.055 ;
        RECT 96.285 215.995 96.575 216.040 ;
        RECT 97.650 215.995 97.970 216.055 ;
        RECT 35.640 215.855 44.980 215.995 ;
        RECT 54.960 215.855 76.720 215.995 ;
        RECT 43.370 215.655 43.690 215.715 ;
        RECT 35.180 215.515 43.690 215.655 ;
        RECT 26.810 215.455 27.130 215.515 ;
        RECT 32.345 215.470 32.635 215.515 ;
        RECT 43.370 215.455 43.690 215.515 ;
        RECT 44.290 215.455 44.610 215.715 ;
        RECT 44.840 215.655 44.980 215.855 ;
        RECT 58.090 215.655 58.410 215.715 ;
        RECT 44.840 215.515 58.410 215.655 ;
        RECT 58.090 215.455 58.410 215.515 ;
        RECT 59.945 215.655 60.235 215.700 ;
        RECT 60.850 215.655 61.170 215.715 ;
        RECT 59.945 215.515 61.170 215.655 ;
        RECT 59.945 215.470 60.235 215.515 ;
        RECT 60.850 215.455 61.170 215.515 ;
        RECT 62.705 215.655 62.995 215.700 ;
        RECT 70.510 215.655 70.830 215.715 ;
        RECT 62.705 215.515 70.830 215.655 ;
        RECT 62.705 215.470 62.995 215.515 ;
        RECT 70.510 215.455 70.830 215.515 ;
        RECT 70.970 215.455 71.290 215.715 ;
        RECT 76.580 215.655 76.720 215.855 ;
        RECT 79.710 215.855 96.040 215.995 ;
        RECT 79.710 215.795 80.030 215.855 ;
        RECT 84.770 215.655 85.090 215.715 ;
        RECT 76.580 215.515 85.090 215.655 ;
        RECT 84.770 215.455 85.090 215.515 ;
        RECT 86.610 215.455 86.930 215.715 ;
        RECT 87.070 215.655 87.390 215.715 ;
        RECT 88.005 215.655 88.295 215.700 ;
        RECT 87.070 215.515 88.295 215.655 ;
        RECT 87.070 215.455 87.390 215.515 ;
        RECT 88.005 215.470 88.295 215.515 ;
        RECT 94.430 215.655 94.750 215.715 ;
        RECT 95.365 215.655 95.655 215.700 ;
        RECT 94.430 215.515 95.655 215.655 ;
        RECT 95.900 215.655 96.040 215.855 ;
        RECT 96.285 215.855 97.970 215.995 ;
        RECT 96.285 215.810 96.575 215.855 ;
        RECT 97.650 215.795 97.970 215.855 ;
        RECT 98.110 215.795 98.430 216.055 ;
        RECT 98.585 215.995 98.875 216.040 ;
        RECT 99.490 215.995 99.810 216.055 ;
        RECT 102.265 215.995 102.555 216.040 ;
        RECT 104.640 215.995 104.780 216.490 ;
        RECT 107.310 216.135 107.630 216.395 ;
        RECT 108.690 216.135 109.010 216.395 ;
        RECT 112.370 216.335 112.690 216.395 ;
        RECT 114.300 216.335 114.440 216.515 ;
        RECT 119.285 216.490 119.575 216.720 ;
        RECT 122.045 216.490 122.335 216.720 ;
        RECT 117.905 216.335 118.195 216.380 ;
        RECT 112.370 216.195 118.195 216.335 ;
        RECT 119.360 216.335 119.500 216.490 ;
        RECT 124.790 216.475 125.110 216.735 ;
        RECT 125.340 216.675 125.480 217.215 ;
        RECT 141.810 217.155 142.130 217.415 ;
        RECT 143.190 217.155 143.510 217.415 ;
        RECT 145.490 217.155 145.810 217.415 ;
        RECT 125.710 217.015 126.030 217.075 ;
        RECT 125.710 216.875 129.620 217.015 ;
        RECT 125.710 216.815 126.030 216.875 ;
        RECT 127.550 216.675 127.870 216.735 ;
        RECT 125.340 216.535 127.870 216.675 ;
        RECT 127.550 216.475 127.870 216.535 ;
        RECT 128.025 216.675 128.315 216.720 ;
        RECT 128.470 216.675 128.790 216.735 ;
        RECT 129.480 216.720 129.620 216.875 ;
        RECT 128.025 216.535 128.790 216.675 ;
        RECT 128.025 216.490 128.315 216.535 ;
        RECT 128.470 216.475 128.790 216.535 ;
        RECT 129.405 216.490 129.695 216.720 ;
        RECT 134.450 216.675 134.770 216.735 ;
        RECT 139.525 216.675 139.815 216.720 ;
        RECT 134.450 216.535 139.815 216.675 ;
        RECT 134.450 216.475 134.770 216.535 ;
        RECT 139.525 216.490 139.815 216.535 ;
        RECT 140.890 216.475 141.210 216.735 ;
        RECT 144.110 216.475 144.430 216.735 ;
        RECT 144.585 216.490 144.875 216.720 ;
        RECT 133.990 216.335 134.310 216.395 ;
        RECT 119.360 216.195 134.310 216.335 ;
        RECT 112.370 216.135 112.690 216.195 ;
        RECT 117.905 216.150 118.195 216.195 ;
        RECT 133.990 216.135 134.310 216.195 ;
        RECT 136.750 216.135 137.070 216.395 ;
        RECT 138.145 216.335 138.435 216.380 ;
        RECT 139.050 216.335 139.370 216.395 ;
        RECT 138.145 216.195 139.370 216.335 ;
        RECT 138.145 216.150 138.435 216.195 ;
        RECT 139.050 216.135 139.370 216.195 ;
        RECT 139.970 216.335 140.290 216.395 ;
        RECT 144.660 216.335 144.800 216.490 ;
        RECT 139.970 216.195 144.800 216.335 ;
        RECT 139.970 216.135 140.290 216.195 ;
        RECT 98.585 215.855 99.810 215.995 ;
        RECT 98.585 215.810 98.875 215.855 ;
        RECT 99.490 215.795 99.810 215.855 ;
        RECT 100.040 215.855 104.780 215.995 ;
        RECT 108.195 215.995 108.485 216.040 ;
        RECT 110.085 215.995 110.375 216.040 ;
        RECT 113.205 215.995 113.495 216.040 ;
        RECT 108.195 215.855 113.495 215.995 ;
        RECT 100.040 215.655 100.180 215.855 ;
        RECT 102.265 215.810 102.555 215.855 ;
        RECT 108.195 215.810 108.485 215.855 ;
        RECT 110.085 215.810 110.375 215.855 ;
        RECT 113.205 215.810 113.495 215.855 ;
        RECT 125.710 215.995 126.030 216.055 ;
        RECT 126.185 215.995 126.475 216.040 ;
        RECT 125.710 215.855 126.475 215.995 ;
        RECT 125.710 215.795 126.030 215.855 ;
        RECT 126.185 215.810 126.475 215.855 ;
        RECT 127.550 215.995 127.870 216.055 ;
        RECT 134.450 215.995 134.770 216.055 ;
        RECT 127.550 215.855 134.770 215.995 ;
        RECT 127.550 215.795 127.870 215.855 ;
        RECT 134.450 215.795 134.770 215.855 ;
        RECT 95.900 215.515 100.180 215.655 ;
        RECT 94.430 215.455 94.750 215.515 ;
        RECT 95.365 215.470 95.655 215.515 ;
        RECT 100.410 215.455 100.730 215.715 ;
        RECT 113.750 215.655 114.070 215.715 ;
        RECT 116.065 215.655 116.355 215.700 ;
        RECT 113.750 215.515 116.355 215.655 ;
        RECT 113.750 215.455 114.070 215.515 ;
        RECT 116.065 215.470 116.355 215.515 ;
        RECT 121.585 215.655 121.875 215.700 ;
        RECT 122.950 215.655 123.270 215.715 ;
        RECT 121.585 215.515 123.270 215.655 ;
        RECT 121.585 215.470 121.875 215.515 ;
        RECT 122.950 215.455 123.270 215.515 ;
        RECT 123.870 215.455 124.190 215.715 ;
        RECT 128.010 215.655 128.330 215.715 ;
        RECT 128.485 215.655 128.775 215.700 ;
        RECT 128.010 215.515 128.775 215.655 ;
        RECT 128.010 215.455 128.330 215.515 ;
        RECT 128.485 215.470 128.775 215.515 ;
        RECT 138.590 215.455 138.910 215.715 ;
        RECT 13.860 214.835 147.720 215.315 ;
        RECT 15.770 214.435 16.090 214.695 ;
        RECT 17.610 214.435 17.930 214.695 ;
        RECT 29.570 214.635 29.890 214.695 ;
        RECT 36.010 214.635 36.330 214.695 ;
        RECT 40.625 214.635 40.915 214.680 ;
        RECT 29.570 214.495 35.780 214.635 ;
        RECT 29.570 214.435 29.890 214.495 ;
        RECT 21.750 214.295 22.070 214.355 ;
        RECT 18.620 214.155 22.070 214.295 ;
        RECT 18.620 213.955 18.760 214.155 ;
        RECT 21.750 214.095 22.070 214.155 ;
        RECT 29.995 214.295 30.285 214.340 ;
        RECT 31.885 214.295 32.175 214.340 ;
        RECT 35.005 214.295 35.295 214.340 ;
        RECT 29.995 214.155 35.295 214.295 ;
        RECT 35.640 214.295 35.780 214.495 ;
        RECT 36.010 214.495 40.915 214.635 ;
        RECT 36.010 214.435 36.330 214.495 ;
        RECT 40.625 214.450 40.915 214.495 ;
        RECT 43.320 214.635 43.610 214.680 ;
        RECT 44.290 214.635 44.610 214.695 ;
        RECT 43.320 214.495 44.610 214.635 ;
        RECT 43.320 214.450 43.610 214.495 ;
        RECT 44.290 214.435 44.610 214.495 ;
        RECT 45.210 214.635 45.530 214.695 ;
        RECT 53.490 214.635 53.810 214.695 ;
        RECT 45.210 214.495 53.810 214.635 ;
        RECT 45.210 214.435 45.530 214.495 ;
        RECT 53.490 214.435 53.810 214.495 ;
        RECT 54.360 214.635 54.650 214.680 ;
        RECT 54.870 214.635 55.190 214.695 ;
        RECT 54.360 214.495 55.190 214.635 ;
        RECT 54.360 214.450 54.650 214.495 ;
        RECT 54.870 214.435 55.190 214.495 ;
        RECT 56.710 214.635 57.030 214.695 ;
        RECT 60.850 214.635 61.170 214.695 ;
        RECT 56.710 214.495 61.170 214.635 ;
        RECT 56.710 214.435 57.030 214.495 ;
        RECT 60.850 214.435 61.170 214.495 ;
        RECT 62.230 214.435 62.550 214.695 ;
        RECT 62.690 214.635 63.010 214.695 ;
        RECT 64.070 214.635 64.390 214.695 ;
        RECT 62.690 214.495 74.420 214.635 ;
        RECT 62.690 214.435 63.010 214.495 ;
        RECT 64.070 214.435 64.390 214.495 ;
        RECT 37.390 214.295 37.710 214.355 ;
        RECT 42.875 214.295 43.165 214.340 ;
        RECT 44.765 214.295 45.055 214.340 ;
        RECT 47.885 214.295 48.175 214.340 ;
        RECT 35.640 214.155 42.680 214.295 ;
        RECT 29.995 214.110 30.285 214.155 ;
        RECT 31.885 214.110 32.175 214.155 ;
        RECT 35.005 214.110 35.295 214.155 ;
        RECT 37.390 214.095 37.710 214.155 ;
        RECT 16.780 213.815 18.760 213.955 ;
        RECT 18.990 213.955 19.310 214.015 ;
        RECT 29.125 213.955 29.415 214.000 ;
        RECT 36.470 213.955 36.790 214.015 ;
        RECT 42.005 213.955 42.295 214.000 ;
        RECT 18.990 213.815 42.295 213.955 ;
        RECT 42.540 213.955 42.680 214.155 ;
        RECT 42.875 214.155 48.175 214.295 ;
        RECT 42.875 214.110 43.165 214.155 ;
        RECT 44.765 214.110 45.055 214.155 ;
        RECT 47.885 214.110 48.175 214.155 ;
        RECT 53.915 214.295 54.205 214.340 ;
        RECT 55.805 214.295 56.095 214.340 ;
        RECT 58.925 214.295 59.215 214.340 ;
        RECT 53.915 214.155 59.215 214.295 ;
        RECT 53.915 214.110 54.205 214.155 ;
        RECT 55.805 214.110 56.095 214.155 ;
        RECT 58.925 214.110 59.215 214.155 ;
        RECT 67.715 214.295 68.005 214.340 ;
        RECT 69.605 214.295 69.895 214.340 ;
        RECT 72.725 214.295 73.015 214.340 ;
        RECT 67.715 214.155 73.015 214.295 ;
        RECT 67.715 214.110 68.005 214.155 ;
        RECT 69.605 214.110 69.895 214.155 ;
        RECT 72.725 214.110 73.015 214.155 ;
        RECT 53.045 213.955 53.335 214.000 ;
        RECT 64.990 213.955 65.310 214.015 ;
        RECT 65.465 213.955 65.755 214.000 ;
        RECT 71.890 213.955 72.210 214.015 ;
        RECT 42.540 213.815 49.580 213.955 ;
        RECT 16.780 213.660 16.920 213.815 ;
        RECT 18.990 213.755 19.310 213.815 ;
        RECT 29.125 213.770 29.415 213.815 ;
        RECT 36.470 213.755 36.790 213.815 ;
        RECT 42.005 213.770 42.295 213.815 ;
        RECT 16.705 213.430 16.995 213.660 ;
        RECT 18.545 213.615 18.835 213.660 ;
        RECT 19.450 213.615 19.770 213.675 ;
        RECT 18.545 213.475 19.770 213.615 ;
        RECT 18.545 213.430 18.835 213.475 ;
        RECT 19.450 213.415 19.770 213.475 ;
        RECT 20.370 213.415 20.690 213.675 ;
        RECT 24.970 213.415 25.290 213.675 ;
        RECT 25.430 213.415 25.750 213.675 ;
        RECT 29.590 213.615 29.880 213.660 ;
        RECT 31.425 213.615 31.715 213.660 ;
        RECT 35.005 213.615 35.295 213.660 ;
        RECT 29.590 213.475 35.295 213.615 ;
        RECT 29.590 213.430 29.880 213.475 ;
        RECT 31.425 213.430 31.715 213.475 ;
        RECT 35.005 213.430 35.295 213.475 ;
        RECT 30.490 213.075 30.810 213.335 ;
        RECT 36.085 213.320 36.375 213.635 ;
        RECT 38.770 213.615 39.090 213.675 ;
        RECT 39.705 213.615 39.995 213.660 ;
        RECT 38.770 213.475 39.995 213.615 ;
        RECT 38.770 213.415 39.090 213.475 ;
        RECT 39.705 213.430 39.995 213.475 ;
        RECT 40.475 213.615 40.765 213.660 ;
        RECT 41.070 213.615 41.390 213.675 ;
        RECT 40.475 213.475 41.390 213.615 ;
        RECT 40.475 213.430 40.765 213.475 ;
        RECT 41.070 213.415 41.390 213.475 ;
        RECT 42.470 213.615 42.760 213.660 ;
        RECT 44.305 213.615 44.595 213.660 ;
        RECT 47.885 213.615 48.175 213.660 ;
        RECT 42.470 213.475 48.175 213.615 ;
        RECT 42.470 213.430 42.760 213.475 ;
        RECT 44.305 213.430 44.595 213.475 ;
        RECT 47.885 213.430 48.175 213.475 ;
        RECT 32.785 213.275 33.435 213.320 ;
        RECT 36.085 213.275 36.675 213.320 ;
        RECT 37.390 213.275 37.710 213.335 ;
        RECT 48.965 213.320 49.255 213.635 ;
        RECT 49.440 213.320 49.580 213.815 ;
        RECT 53.045 213.815 64.300 213.955 ;
        RECT 53.045 213.770 53.335 213.815 ;
        RECT 53.510 213.615 53.800 213.660 ;
        RECT 55.345 213.615 55.635 213.660 ;
        RECT 58.925 213.615 59.215 213.660 ;
        RECT 53.510 213.475 59.215 213.615 ;
        RECT 53.510 213.430 53.800 213.475 ;
        RECT 55.345 213.430 55.635 213.475 ;
        RECT 58.925 213.430 59.215 213.475 ;
        RECT 60.005 213.615 60.295 213.635 ;
        RECT 60.850 213.615 61.170 213.675 ;
        RECT 63.610 213.615 63.930 213.675 ;
        RECT 60.005 213.475 63.930 213.615 ;
        RECT 64.160 213.615 64.300 213.815 ;
        RECT 64.990 213.815 72.210 213.955 ;
        RECT 64.990 213.755 65.310 213.815 ;
        RECT 65.465 213.770 65.755 213.815 ;
        RECT 71.890 213.755 72.210 213.815 ;
        RECT 66.830 213.615 67.150 213.675 ;
        RECT 64.160 213.475 67.150 213.615 ;
        RECT 56.710 213.320 57.030 213.335 ;
        RECT 60.005 213.320 60.295 213.475 ;
        RECT 60.850 213.415 61.170 213.475 ;
        RECT 63.610 213.415 63.930 213.475 ;
        RECT 66.830 213.415 67.150 213.475 ;
        RECT 67.310 213.615 67.600 213.660 ;
        RECT 69.145 213.615 69.435 213.660 ;
        RECT 72.725 213.615 73.015 213.660 ;
        RECT 67.310 213.475 73.015 213.615 ;
        RECT 67.310 213.430 67.600 213.475 ;
        RECT 69.145 213.430 69.435 213.475 ;
        RECT 72.725 213.430 73.015 213.475 ;
        RECT 32.785 213.135 37.710 213.275 ;
        RECT 32.785 213.090 33.435 213.135 ;
        RECT 36.385 213.090 36.675 213.135 ;
        RECT 37.390 213.075 37.710 213.135 ;
        RECT 39.245 213.090 39.535 213.320 ;
        RECT 45.665 213.275 46.315 213.320 ;
        RECT 48.965 213.275 49.580 213.320 ;
        RECT 56.705 213.275 57.355 213.320 ;
        RECT 60.005 213.275 60.595 213.320 ;
        RECT 64.085 213.275 64.375 213.320 ;
        RECT 45.665 213.135 60.595 213.275 ;
        RECT 45.665 213.090 46.315 213.135 ;
        RECT 49.265 213.090 49.555 213.135 ;
        RECT 56.705 213.090 57.355 213.135 ;
        RECT 60.305 213.090 60.595 213.135 ;
        RECT 60.940 213.135 62.460 213.275 ;
        RECT 14.390 212.935 14.710 212.995 ;
        RECT 19.465 212.935 19.755 212.980 ;
        RECT 14.390 212.795 19.755 212.935 ;
        RECT 14.390 212.735 14.710 212.795 ;
        RECT 19.465 212.750 19.755 212.795 ;
        RECT 26.365 212.935 26.655 212.980 ;
        RECT 36.930 212.935 37.250 212.995 ;
        RECT 26.365 212.795 37.250 212.935 ;
        RECT 39.320 212.935 39.460 213.090 ;
        RECT 56.710 213.075 57.030 213.090 ;
        RECT 39.690 212.935 40.010 212.995 ;
        RECT 39.320 212.795 40.010 212.935 ;
        RECT 26.365 212.750 26.655 212.795 ;
        RECT 36.930 212.735 37.250 212.795 ;
        RECT 39.690 212.735 40.010 212.795 ;
        RECT 49.810 212.935 50.130 212.995 ;
        RECT 50.745 212.935 51.035 212.980 ;
        RECT 60.940 212.935 61.080 213.135 ;
        RECT 49.810 212.795 61.080 212.935 ;
        RECT 61.310 212.935 61.630 212.995 ;
        RECT 61.785 212.935 62.075 212.980 ;
        RECT 61.310 212.795 62.075 212.935 ;
        RECT 62.320 212.935 62.460 213.135 ;
        RECT 64.085 213.135 67.980 213.275 ;
        RECT 64.085 213.090 64.375 213.135 ;
        RECT 64.545 212.935 64.835 212.980 ;
        RECT 62.320 212.795 64.835 212.935 ;
        RECT 67.840 212.935 67.980 213.135 ;
        RECT 68.210 213.075 68.530 213.335 ;
        RECT 73.805 213.320 74.095 213.635 ;
        RECT 74.280 213.320 74.420 214.495 ;
        RECT 79.250 214.435 79.570 214.695 ;
        RECT 81.090 214.635 81.410 214.695 ;
        RECT 86.685 214.635 86.975 214.680 ;
        RECT 81.090 214.495 86.975 214.635 ;
        RECT 81.090 214.435 81.410 214.495 ;
        RECT 86.685 214.450 86.975 214.495 ;
        RECT 97.190 214.435 97.510 214.695 ;
        RECT 99.505 214.635 99.795 214.680 ;
        RECT 108.690 214.635 109.010 214.695 ;
        RECT 111.005 214.635 111.295 214.680 ;
        RECT 99.505 214.495 102.020 214.635 ;
        RECT 99.505 214.450 99.795 214.495 ;
        RECT 82.125 214.295 82.415 214.340 ;
        RECT 85.245 214.295 85.535 214.340 ;
        RECT 87.135 214.295 87.425 214.340 ;
        RECT 82.125 214.155 87.425 214.295 ;
        RECT 82.125 214.110 82.415 214.155 ;
        RECT 85.245 214.110 85.535 214.155 ;
        RECT 87.135 214.110 87.425 214.155 ;
        RECT 89.335 214.295 89.625 214.340 ;
        RECT 91.225 214.295 91.515 214.340 ;
        RECT 94.345 214.295 94.635 214.340 ;
        RECT 89.335 214.155 94.635 214.295 ;
        RECT 89.335 214.110 89.625 214.155 ;
        RECT 91.225 214.110 91.515 214.155 ;
        RECT 94.345 214.110 94.635 214.155 ;
        RECT 74.650 213.955 74.970 214.015 ;
        RECT 76.965 213.955 77.255 214.000 ;
        RECT 74.650 213.815 77.255 213.955 ;
        RECT 74.650 213.755 74.970 213.815 ;
        RECT 76.965 213.770 77.255 213.815 ;
        RECT 86.150 213.955 86.470 214.015 ;
        RECT 97.280 213.955 97.420 214.435 ;
        RECT 99.950 214.095 100.270 214.355 ;
        RECT 101.330 213.955 101.650 214.015 ;
        RECT 86.150 213.815 96.040 213.955 ;
        RECT 97.280 213.815 101.650 213.955 ;
        RECT 101.880 213.955 102.020 214.495 ;
        RECT 108.690 214.495 111.295 214.635 ;
        RECT 108.690 214.435 109.010 214.495 ;
        RECT 111.005 214.450 111.295 214.495 ;
        RECT 119.725 214.635 120.015 214.680 ;
        RECT 120.645 214.635 120.935 214.680 ;
        RECT 119.725 214.495 120.935 214.635 ;
        RECT 119.725 214.450 120.015 214.495 ;
        RECT 120.645 214.450 120.935 214.495 ;
        RECT 121.570 214.635 121.890 214.695 ;
        RECT 139.970 214.635 140.290 214.695 ;
        RECT 121.570 214.495 140.290 214.635 ;
        RECT 121.570 214.435 121.890 214.495 ;
        RECT 139.970 214.435 140.290 214.495 ;
        RECT 102.710 214.295 103.030 214.355 ;
        RECT 131.195 214.295 131.485 214.340 ;
        RECT 133.085 214.295 133.375 214.340 ;
        RECT 136.205 214.295 136.495 214.340 ;
        RECT 102.710 214.155 105.240 214.295 ;
        RECT 102.710 214.095 103.030 214.155 ;
        RECT 102.265 213.955 102.555 214.000 ;
        RECT 101.880 213.815 102.555 213.955 ;
        RECT 86.150 213.755 86.470 213.815 ;
        RECT 75.110 213.615 75.430 213.675 ;
        RECT 76.505 213.615 76.795 213.660 ;
        RECT 75.110 213.475 76.795 213.615 ;
        RECT 75.110 213.415 75.430 213.475 ;
        RECT 76.505 213.430 76.795 213.475 ;
        RECT 70.505 213.275 71.155 213.320 ;
        RECT 73.805 213.275 74.420 213.320 ;
        RECT 79.710 213.275 80.030 213.335 ;
        RECT 81.045 213.320 81.335 213.635 ;
        RECT 82.125 213.615 82.415 213.660 ;
        RECT 85.705 213.615 85.995 213.660 ;
        RECT 87.540 213.615 87.830 213.660 ;
        RECT 82.125 213.475 87.830 213.615 ;
        RECT 82.125 213.430 82.415 213.475 ;
        RECT 85.705 213.430 85.995 213.475 ;
        RECT 87.540 213.430 87.830 213.475 ;
        RECT 88.005 213.615 88.295 213.660 ;
        RECT 88.450 213.615 88.770 213.675 ;
        RECT 88.005 213.475 88.770 213.615 ;
        RECT 88.005 213.430 88.295 213.475 ;
        RECT 88.450 213.415 88.770 213.475 ;
        RECT 88.930 213.615 89.220 213.660 ;
        RECT 90.765 213.615 91.055 213.660 ;
        RECT 94.345 213.615 94.635 213.660 ;
        RECT 88.930 213.475 94.635 213.615 ;
        RECT 88.930 213.430 89.220 213.475 ;
        RECT 90.765 213.430 91.055 213.475 ;
        RECT 94.345 213.430 94.635 213.475 ;
        RECT 70.505 213.135 80.030 213.275 ;
        RECT 70.505 213.090 71.155 213.135 ;
        RECT 74.105 213.090 74.395 213.135 ;
        RECT 79.710 213.075 80.030 213.135 ;
        RECT 80.745 213.275 81.335 213.320 ;
        RECT 83.985 213.275 84.635 213.320 ;
        RECT 85.230 213.275 85.550 213.335 ;
        RECT 80.745 213.135 89.600 213.275 ;
        RECT 80.745 213.090 81.035 213.135 ;
        RECT 83.985 213.090 84.635 213.135 ;
        RECT 85.230 213.075 85.550 213.135 ;
        RECT 72.350 212.935 72.670 212.995 ;
        RECT 67.840 212.795 72.670 212.935 ;
        RECT 49.810 212.735 50.130 212.795 ;
        RECT 50.745 212.750 51.035 212.795 ;
        RECT 61.310 212.735 61.630 212.795 ;
        RECT 61.785 212.750 62.075 212.795 ;
        RECT 64.545 212.750 64.835 212.795 ;
        RECT 72.350 212.735 72.670 212.795 ;
        RECT 75.110 212.935 75.430 212.995 ;
        RECT 75.585 212.935 75.875 212.980 ;
        RECT 75.110 212.795 75.875 212.935 ;
        RECT 89.460 212.935 89.600 213.135 ;
        RECT 89.830 213.075 90.150 213.335 ;
        RECT 95.425 213.320 95.715 213.635 ;
        RECT 95.900 213.615 96.040 213.815 ;
        RECT 101.330 213.755 101.650 213.815 ;
        RECT 102.265 213.770 102.555 213.815 ;
        RECT 103.185 213.955 103.475 214.000 ;
        RECT 104.565 213.955 104.855 214.000 ;
        RECT 103.185 213.815 104.855 213.955 ;
        RECT 105.100 213.955 105.240 214.155 ;
        RECT 131.195 214.155 136.495 214.295 ;
        RECT 131.195 214.110 131.485 214.155 ;
        RECT 133.085 214.110 133.375 214.155 ;
        RECT 136.205 214.110 136.495 214.155 ;
        RECT 105.100 213.815 107.540 213.955 ;
        RECT 103.185 213.770 103.475 213.815 ;
        RECT 104.565 213.770 104.855 213.815 ;
        RECT 97.665 213.615 97.955 213.660 ;
        RECT 95.900 213.475 97.955 213.615 ;
        RECT 97.665 213.430 97.955 213.475 ;
        RECT 98.585 213.615 98.875 213.660 ;
        RECT 100.870 213.615 101.190 213.675 ;
        RECT 98.585 213.475 101.190 213.615 ;
        RECT 98.585 213.430 98.875 213.475 ;
        RECT 92.125 213.275 92.775 213.320 ;
        RECT 95.425 213.275 96.015 213.320 ;
        RECT 97.740 213.275 97.880 213.430 ;
        RECT 100.870 213.415 101.190 213.475 ;
        RECT 101.790 213.415 102.110 213.675 ;
        RECT 105.485 213.615 105.775 213.660 ;
        RECT 106.390 213.615 106.710 213.675 ;
        RECT 105.485 213.475 106.710 213.615 ;
        RECT 105.485 213.430 105.775 213.475 ;
        RECT 106.390 213.415 106.710 213.475 ;
        RECT 106.850 213.415 107.170 213.675 ;
        RECT 107.400 213.615 107.540 213.815 ;
        RECT 114.210 213.755 114.530 214.015 ;
        RECT 117.430 213.755 117.750 214.015 ;
        RECT 120.190 213.755 120.510 214.015 ;
        RECT 122.030 213.955 122.350 214.015 ;
        RECT 127.550 213.955 127.870 214.015 ;
        RECT 122.030 213.815 127.870 213.955 ;
        RECT 122.030 213.755 122.350 213.815 ;
        RECT 108.690 213.615 109.010 213.675 ;
        RECT 124.880 213.660 125.020 213.815 ;
        RECT 127.550 213.755 127.870 213.815 ;
        RECT 131.690 213.955 132.010 214.015 ;
        RECT 146.410 213.955 146.730 214.015 ;
        RECT 131.690 213.815 142.040 213.955 ;
        RECT 131.690 213.755 132.010 213.815 ;
        RECT 116.065 213.615 116.355 213.660 ;
        RECT 121.585 213.615 121.875 213.660 ;
        RECT 107.400 213.475 121.875 213.615 ;
        RECT 108.690 213.415 109.010 213.475 ;
        RECT 116.065 213.430 116.355 213.475 ;
        RECT 121.585 213.430 121.875 213.475 ;
        RECT 124.800 213.430 125.090 213.660 ;
        RECT 125.265 213.430 125.555 213.660 ;
        RECT 104.090 213.275 104.410 213.335 ;
        RECT 107.325 213.275 107.615 213.320 ;
        RECT 92.125 213.135 97.420 213.275 ;
        RECT 97.740 213.135 98.800 213.275 ;
        RECT 92.125 213.090 92.775 213.135 ;
        RECT 95.725 213.090 96.015 213.135 ;
        RECT 97.280 212.935 97.420 213.135 ;
        RECT 98.110 212.935 98.430 212.995 ;
        RECT 89.460 212.795 98.430 212.935 ;
        RECT 98.660 212.935 98.800 213.135 ;
        RECT 104.090 213.135 107.615 213.275 ;
        RECT 104.090 213.075 104.410 213.135 ;
        RECT 107.325 213.090 107.615 213.135 ;
        RECT 108.230 213.075 108.550 213.335 ;
        RECT 116.525 213.275 116.815 213.320 ;
        RECT 120.190 213.275 120.510 213.335 ;
        RECT 116.525 213.135 120.510 213.275 ;
        RECT 121.660 213.275 121.800 213.430 ;
        RECT 122.950 213.275 123.270 213.335 ;
        RECT 121.660 213.135 123.270 213.275 ;
        RECT 116.525 213.090 116.815 213.135 ;
        RECT 120.190 213.075 120.510 213.135 ;
        RECT 122.950 213.075 123.270 213.135 ;
        RECT 123.870 213.275 124.190 213.335 ;
        RECT 125.340 213.275 125.480 213.430 ;
        RECT 127.090 213.415 127.410 213.675 ;
        RECT 128.010 213.415 128.330 213.675 ;
        RECT 128.485 213.430 128.775 213.660 ;
        RECT 123.870 213.135 125.480 213.275 ;
        RECT 123.870 213.075 124.190 213.135 ;
        RECT 105.010 212.935 105.330 212.995 ;
        RECT 98.660 212.795 105.330 212.935 ;
        RECT 75.110 212.735 75.430 212.795 ;
        RECT 75.585 212.750 75.875 212.795 ;
        RECT 98.110 212.735 98.430 212.795 ;
        RECT 105.010 212.735 105.330 212.795 ;
        RECT 105.930 212.935 106.250 212.995 ;
        RECT 106.405 212.935 106.695 212.980 ;
        RECT 105.930 212.795 106.695 212.935 ;
        RECT 105.930 212.735 106.250 212.795 ;
        RECT 106.405 212.750 106.695 212.795 ;
        RECT 112.830 212.735 113.150 212.995 ;
        RECT 113.290 212.735 113.610 212.995 ;
        RECT 121.110 212.935 121.430 212.995 ;
        RECT 123.425 212.935 123.715 212.980 ;
        RECT 121.110 212.795 123.715 212.935 ;
        RECT 121.110 212.735 121.430 212.795 ;
        RECT 123.425 212.750 123.715 212.795 ;
        RECT 125.250 212.935 125.570 212.995 ;
        RECT 126.185 212.935 126.475 212.980 ;
        RECT 125.250 212.795 126.475 212.935 ;
        RECT 128.560 212.935 128.700 213.430 ;
        RECT 130.310 213.415 130.630 213.675 ;
        RECT 130.790 213.615 131.080 213.660 ;
        RECT 132.625 213.615 132.915 213.660 ;
        RECT 136.205 213.615 136.495 213.660 ;
        RECT 130.790 213.475 136.495 213.615 ;
        RECT 130.790 213.430 131.080 213.475 ;
        RECT 132.625 213.430 132.915 213.475 ;
        RECT 136.205 213.430 136.495 213.475 ;
        RECT 131.705 213.275 131.995 213.320 ;
        RECT 133.070 213.275 133.390 213.335 ;
        RECT 133.990 213.320 134.310 213.335 ;
        RECT 137.285 213.320 137.575 213.635 ;
        RECT 140.890 213.415 141.210 213.675 ;
        RECT 131.705 213.135 133.390 213.275 ;
        RECT 131.705 213.090 131.995 213.135 ;
        RECT 133.070 213.075 133.390 213.135 ;
        RECT 133.985 213.275 134.635 213.320 ;
        RECT 137.285 213.275 137.875 213.320 ;
        RECT 133.985 213.135 137.875 213.275 ;
        RECT 133.985 213.090 134.635 213.135 ;
        RECT 137.585 213.090 137.875 213.135 ;
        RECT 138.130 213.275 138.450 213.335 ;
        RECT 141.900 213.275 142.040 213.815 ;
        RECT 142.360 213.815 146.730 213.955 ;
        RECT 142.360 213.660 142.500 213.815 ;
        RECT 146.410 213.755 146.730 213.815 ;
        RECT 142.285 213.430 142.575 213.660 ;
        RECT 142.730 213.415 143.050 213.675 ;
        RECT 144.585 213.430 144.875 213.660 ;
        RECT 144.660 213.275 144.800 213.430 ;
        RECT 138.130 213.135 141.580 213.275 ;
        RECT 141.900 213.135 144.800 213.275 ;
        RECT 133.990 213.075 134.310 213.090 ;
        RECT 138.130 213.075 138.450 213.135 ;
        RECT 135.830 212.935 136.150 212.995 ;
        RECT 128.560 212.795 136.150 212.935 ;
        RECT 125.250 212.735 125.570 212.795 ;
        RECT 126.185 212.750 126.475 212.795 ;
        RECT 135.830 212.735 136.150 212.795 ;
        RECT 139.050 212.735 139.370 212.995 ;
        RECT 139.970 212.735 140.290 212.995 ;
        RECT 141.440 212.980 141.580 213.135 ;
        RECT 141.365 212.750 141.655 212.980 ;
        RECT 143.650 212.735 143.970 212.995 ;
        RECT 145.505 212.935 145.795 212.980 ;
        RECT 145.950 212.935 146.270 212.995 ;
        RECT 145.505 212.795 146.270 212.935 ;
        RECT 145.505 212.750 145.795 212.795 ;
        RECT 145.950 212.735 146.270 212.795 ;
        RECT 13.860 212.115 147.720 212.595 ;
        RECT 14.850 211.915 15.170 211.975 ;
        RECT 15.785 211.915 16.075 211.960 ;
        RECT 30.490 211.915 30.810 211.975 ;
        RECT 31.425 211.915 31.715 211.960 ;
        RECT 14.850 211.775 16.075 211.915 ;
        RECT 14.850 211.715 15.170 211.775 ;
        RECT 15.785 211.730 16.075 211.775 ;
        RECT 18.160 211.775 30.260 211.915 ;
        RECT 16.705 211.235 16.995 211.280 ;
        RECT 18.160 211.235 18.300 211.775 ;
        RECT 22.665 211.575 23.315 211.620 ;
        RECT 26.265 211.575 26.555 211.620 ;
        RECT 29.570 211.575 29.890 211.635 ;
        RECT 22.665 211.435 29.890 211.575 ;
        RECT 30.120 211.575 30.260 211.775 ;
        RECT 30.490 211.775 31.715 211.915 ;
        RECT 30.490 211.715 30.810 211.775 ;
        RECT 31.425 211.730 31.715 211.775 ;
        RECT 33.250 211.915 33.570 211.975 ;
        RECT 36.930 211.915 37.250 211.975 ;
        RECT 33.250 211.775 37.250 211.915 ;
        RECT 33.250 211.715 33.570 211.775 ;
        RECT 36.930 211.715 37.250 211.775 ;
        RECT 46.590 211.915 46.910 211.975 ;
        RECT 47.985 211.915 48.275 211.960 ;
        RECT 46.590 211.775 48.275 211.915 ;
        RECT 46.590 211.715 46.910 211.775 ;
        RECT 47.985 211.730 48.275 211.775 ;
        RECT 48.890 211.915 49.210 211.975 ;
        RECT 48.890 211.775 52.340 211.915 ;
        RECT 48.890 211.715 49.210 211.775 ;
        RECT 36.010 211.575 36.330 211.635 ;
        RECT 30.120 211.435 36.330 211.575 ;
        RECT 22.665 211.390 23.315 211.435 ;
        RECT 25.965 211.390 26.555 211.435 ;
        RECT 16.705 211.095 18.300 211.235 ;
        RECT 16.705 211.050 16.995 211.095 ;
        RECT 18.530 211.035 18.850 211.295 ;
        RECT 18.990 211.035 19.310 211.295 ;
        RECT 19.470 211.235 19.760 211.280 ;
        RECT 21.305 211.235 21.595 211.280 ;
        RECT 24.885 211.235 25.175 211.280 ;
        RECT 19.470 211.095 25.175 211.235 ;
        RECT 19.470 211.050 19.760 211.095 ;
        RECT 21.305 211.050 21.595 211.095 ;
        RECT 24.885 211.050 25.175 211.095 ;
        RECT 25.965 211.075 26.255 211.390 ;
        RECT 20.385 210.895 20.675 210.940 ;
        RECT 27.270 210.895 27.590 210.955 ;
        RECT 20.385 210.755 27.590 210.895 ;
        RECT 20.385 210.710 20.675 210.755 ;
        RECT 27.270 210.695 27.590 210.755 ;
        RECT 14.510 210.555 14.830 210.615 ;
        RECT 17.625 210.555 17.915 210.600 ;
        RECT 14.510 210.415 17.915 210.555 ;
        RECT 14.510 210.355 14.830 210.415 ;
        RECT 17.625 210.370 17.915 210.415 ;
        RECT 19.875 210.555 20.165 210.600 ;
        RECT 21.765 210.555 22.055 210.600 ;
        RECT 24.885 210.555 25.175 210.600 ;
        RECT 19.875 210.415 25.175 210.555 ;
        RECT 19.875 210.370 20.165 210.415 ;
        RECT 21.765 210.370 22.055 210.415 ;
        RECT 24.885 210.370 25.175 210.415 ;
        RECT 26.350 210.555 26.670 210.615 ;
        RECT 27.820 210.555 27.960 211.435 ;
        RECT 29.570 211.375 29.890 211.435 ;
        RECT 36.010 211.375 36.330 211.435 ;
        RECT 47.065 211.575 47.355 211.620 ;
        RECT 51.650 211.575 51.970 211.635 ;
        RECT 47.065 211.435 51.970 211.575 ;
        RECT 52.200 211.575 52.340 211.775 ;
        RECT 54.870 211.715 55.190 211.975 ;
        RECT 56.710 211.915 57.030 211.975 ;
        RECT 56.570 211.715 57.030 211.915 ;
        RECT 61.310 211.915 61.630 211.975 ;
        RECT 61.785 211.915 62.075 211.960 ;
        RECT 61.310 211.775 62.075 211.915 ;
        RECT 61.310 211.715 61.630 211.775 ;
        RECT 61.785 211.730 62.075 211.775 ;
        RECT 62.230 211.715 62.550 211.975 ;
        RECT 64.085 211.915 64.375 211.960 ;
        RECT 64.530 211.915 64.850 211.975 ;
        RECT 64.085 211.775 64.850 211.915 ;
        RECT 64.085 211.730 64.375 211.775 ;
        RECT 64.530 211.715 64.850 211.775 ;
        RECT 68.210 211.915 68.530 211.975 ;
        RECT 69.145 211.915 69.435 211.960 ;
        RECT 68.210 211.775 69.435 211.915 ;
        RECT 68.210 211.715 68.530 211.775 ;
        RECT 69.145 211.730 69.435 211.775 ;
        RECT 70.970 211.915 71.290 211.975 ;
        RECT 71.445 211.915 71.735 211.960 ;
        RECT 70.970 211.775 71.735 211.915 ;
        RECT 70.970 211.715 71.290 211.775 ;
        RECT 71.445 211.730 71.735 211.775 ;
        RECT 78.790 211.915 79.110 211.975 ;
        RECT 79.265 211.915 79.555 211.960 ;
        RECT 78.790 211.775 79.555 211.915 ;
        RECT 78.790 211.715 79.110 211.775 ;
        RECT 79.265 211.730 79.555 211.775 ;
        RECT 81.090 211.715 81.410 211.975 ;
        RECT 82.470 211.915 82.790 211.975 ;
        RECT 85.230 211.915 85.550 211.975 ;
        RECT 82.470 211.775 85.550 211.915 ;
        RECT 82.470 211.715 82.790 211.775 ;
        RECT 85.230 211.715 85.550 211.775 ;
        RECT 86.610 211.915 86.930 211.975 ;
        RECT 87.085 211.915 87.375 211.960 ;
        RECT 86.610 211.775 87.375 211.915 ;
        RECT 86.610 211.715 86.930 211.775 ;
        RECT 87.085 211.730 87.375 211.775 ;
        RECT 88.925 211.915 89.215 211.960 ;
        RECT 89.830 211.915 90.150 211.975 ;
        RECT 98.570 211.915 98.890 211.975 ;
        RECT 104.090 211.915 104.410 211.975 ;
        RECT 88.925 211.775 90.150 211.915 ;
        RECT 88.925 211.730 89.215 211.775 ;
        RECT 89.830 211.715 90.150 211.775 ;
        RECT 97.740 211.775 104.410 211.915 ;
        RECT 56.570 211.575 56.710 211.715 ;
        RECT 52.200 211.435 56.710 211.575 ;
        RECT 57.170 211.575 57.490 211.635 ;
        RECT 60.850 211.575 61.170 211.635 ;
        RECT 65.910 211.575 66.230 211.635 ;
        RECT 57.170 211.435 66.230 211.575 ;
        RECT 47.065 211.390 47.355 211.435 ;
        RECT 51.650 211.375 51.970 211.435 ;
        RECT 57.170 211.375 57.490 211.435 ;
        RECT 35.090 211.235 35.410 211.295 ;
        RECT 36.485 211.235 36.775 211.280 ;
        RECT 35.090 211.095 36.775 211.235 ;
        RECT 35.090 211.035 35.410 211.095 ;
        RECT 36.485 211.050 36.775 211.095 ;
        RECT 37.850 211.035 38.170 211.295 ;
        RECT 48.890 211.235 49.210 211.295 ;
        RECT 38.860 211.095 49.210 211.235 ;
        RECT 29.125 210.895 29.415 210.940 ;
        RECT 32.330 210.895 32.650 210.955 ;
        RECT 29.125 210.755 32.650 210.895 ;
        RECT 29.125 210.710 29.415 210.755 ;
        RECT 32.330 210.695 32.650 210.755 ;
        RECT 33.725 210.710 34.015 210.940 ;
        RECT 34.645 210.895 34.935 210.940 ;
        RECT 35.565 210.895 35.855 210.940 ;
        RECT 34.645 210.755 35.855 210.895 ;
        RECT 34.645 210.710 34.935 210.755 ;
        RECT 35.565 210.710 35.855 210.755 ;
        RECT 36.010 210.895 36.330 210.955 ;
        RECT 36.945 210.895 37.235 210.940 ;
        RECT 36.010 210.755 37.235 210.895 ;
        RECT 26.350 210.415 27.960 210.555 ;
        RECT 31.870 210.555 32.190 210.615 ;
        RECT 33.800 210.555 33.940 210.710 ;
        RECT 36.010 210.695 36.330 210.755 ;
        RECT 36.945 210.710 37.235 210.755 ;
        RECT 37.390 210.895 37.710 210.955 ;
        RECT 38.860 210.895 39.000 211.095 ;
        RECT 48.890 211.035 49.210 211.095 ;
        RECT 49.810 211.035 50.130 211.295 ;
        RECT 50.730 211.235 51.050 211.295 ;
        RECT 51.205 211.235 51.495 211.280 ;
        RECT 50.730 211.095 51.495 211.235 ;
        RECT 50.730 211.035 51.050 211.095 ;
        RECT 51.205 211.050 51.495 211.095 ;
        RECT 52.110 211.035 52.430 211.295 ;
        RECT 54.425 211.050 54.715 211.280 ;
        RECT 55.330 211.235 55.650 211.295 ;
        RECT 60.020 211.280 60.160 211.435 ;
        RECT 60.850 211.375 61.170 211.435 ;
        RECT 65.910 211.375 66.230 211.435 ;
        RECT 69.590 211.575 69.910 211.635 ;
        RECT 75.110 211.575 75.430 211.635 ;
        RECT 91.210 211.575 91.530 211.635 ;
        RECT 92.145 211.575 92.435 211.620 ;
        RECT 96.730 211.575 97.050 211.635 ;
        RECT 69.590 211.435 75.430 211.575 ;
        RECT 69.590 211.375 69.910 211.435 ;
        RECT 56.725 211.235 57.015 211.280 ;
        RECT 55.330 211.095 59.700 211.235 ;
        RECT 37.390 210.755 39.000 210.895 ;
        RECT 40.150 210.895 40.470 210.955 ;
        RECT 40.625 210.895 40.915 210.940 ;
        RECT 40.150 210.755 40.915 210.895 ;
        RECT 37.390 210.695 37.710 210.755 ;
        RECT 40.150 210.695 40.470 210.755 ;
        RECT 40.625 210.710 40.915 210.755 ;
        RECT 41.990 210.695 42.310 210.955 ;
        RECT 54.500 210.895 54.640 211.050 ;
        RECT 55.330 211.035 55.650 211.095 ;
        RECT 56.725 211.050 57.015 211.095 ;
        RECT 54.870 210.895 55.190 210.955 ;
        RECT 54.500 210.755 55.190 210.895 ;
        RECT 54.870 210.695 55.190 210.755 ;
        RECT 55.790 210.895 56.110 210.955 ;
        RECT 57.185 210.895 57.475 210.940 ;
        RECT 55.790 210.755 57.475 210.895 ;
        RECT 55.790 210.695 56.110 210.755 ;
        RECT 57.185 210.710 57.475 210.755 ;
        RECT 57.630 210.695 57.950 210.955 ;
        RECT 59.560 210.895 59.700 211.095 ;
        RECT 59.945 211.050 60.235 211.280 ;
        RECT 67.750 211.235 68.070 211.295 ;
        RECT 70.985 211.235 71.275 211.280 ;
        RECT 73.285 211.235 73.575 211.280 ;
        RECT 73.730 211.235 74.050 211.295 ;
        RECT 60.480 211.095 73.040 211.235 ;
        RECT 60.480 210.895 60.620 211.095 ;
        RECT 67.750 211.035 68.070 211.095 ;
        RECT 70.985 211.050 71.275 211.095 ;
        RECT 59.560 210.755 60.620 210.895 ;
        RECT 60.850 210.695 61.170 210.955 ;
        RECT 63.150 210.895 63.470 210.955 ;
        RECT 70.050 210.895 70.370 210.955 ;
        RECT 63.150 210.755 70.370 210.895 ;
        RECT 63.150 210.695 63.470 210.755 ;
        RECT 70.050 210.695 70.370 210.755 ;
        RECT 72.365 210.710 72.655 210.940 ;
        RECT 72.900 210.895 73.040 211.095 ;
        RECT 73.285 211.095 74.050 211.235 ;
        RECT 73.285 211.050 73.575 211.095 ;
        RECT 73.730 211.035 74.050 211.095 ;
        RECT 74.190 211.035 74.510 211.295 ;
        RECT 74.740 211.235 74.880 211.435 ;
        RECT 75.110 211.375 75.430 211.435 ;
        RECT 76.120 211.435 86.840 211.575 ;
        RECT 75.585 211.235 75.875 211.280 ;
        RECT 74.740 211.095 75.875 211.235 ;
        RECT 75.585 211.050 75.875 211.095 ;
        RECT 76.120 210.895 76.260 211.435 ;
        RECT 76.490 211.035 76.810 211.295 ;
        RECT 82.010 211.035 82.330 211.295 ;
        RECT 84.325 211.235 84.615 211.280 ;
        RECT 84.770 211.235 85.090 211.295 ;
        RECT 86.700 211.280 86.840 211.435 ;
        RECT 91.210 211.435 92.435 211.575 ;
        RECT 91.210 211.375 91.530 211.435 ;
        RECT 92.145 211.390 92.435 211.435 ;
        RECT 94.520 211.435 97.050 211.575 ;
        RECT 94.520 211.295 94.660 211.435 ;
        RECT 96.730 211.375 97.050 211.435 ;
        RECT 97.190 211.375 97.510 211.635 ;
        RECT 84.325 211.095 85.090 211.235 ;
        RECT 84.325 211.050 84.615 211.095 ;
        RECT 84.770 211.035 85.090 211.095 ;
        RECT 86.625 211.235 86.915 211.280 ;
        RECT 87.070 211.235 87.390 211.295 ;
        RECT 86.625 211.095 87.390 211.235 ;
        RECT 86.625 211.050 86.915 211.095 ;
        RECT 87.070 211.035 87.390 211.095 ;
        RECT 87.530 211.235 87.850 211.295 ;
        RECT 89.385 211.235 89.675 211.280 ;
        RECT 87.530 211.095 89.675 211.235 ;
        RECT 87.530 211.035 87.850 211.095 ;
        RECT 89.385 211.050 89.675 211.095 ;
        RECT 90.305 211.235 90.595 211.280 ;
        RECT 90.750 211.235 91.070 211.295 ;
        RECT 90.305 211.095 91.070 211.235 ;
        RECT 90.305 211.050 90.595 211.095 ;
        RECT 90.750 211.035 91.070 211.095 ;
        RECT 93.050 211.035 93.370 211.295 ;
        RECT 94.430 211.035 94.750 211.295 ;
        RECT 95.825 211.235 96.115 211.280 ;
        RECT 97.740 211.235 97.880 211.775 ;
        RECT 98.570 211.715 98.890 211.775 ;
        RECT 104.090 211.715 104.410 211.775 ;
        RECT 105.010 211.915 105.330 211.975 ;
        RECT 107.325 211.915 107.615 211.960 ;
        RECT 109.610 211.915 109.930 211.975 ;
        RECT 105.010 211.775 109.930 211.915 ;
        RECT 105.010 211.715 105.330 211.775 ;
        RECT 107.325 211.730 107.615 211.775 ;
        RECT 109.610 211.715 109.930 211.775 ;
        RECT 114.210 211.915 114.530 211.975 ;
        RECT 122.045 211.915 122.335 211.960 ;
        RECT 124.790 211.915 125.110 211.975 ;
        RECT 132.610 211.915 132.930 211.975 ;
        RECT 114.210 211.775 122.335 211.915 ;
        RECT 114.210 211.715 114.530 211.775 ;
        RECT 122.045 211.730 122.335 211.775 ;
        RECT 123.500 211.775 132.930 211.915 ;
        RECT 99.950 211.375 100.270 211.635 ;
        RECT 102.245 211.575 102.895 211.620 ;
        RECT 105.845 211.575 106.135 211.620 ;
        RECT 122.490 211.575 122.810 211.635 ;
        RECT 102.245 211.435 106.135 211.575 ;
        RECT 102.245 211.390 102.895 211.435 ;
        RECT 105.545 211.390 106.135 211.435 ;
        RECT 120.740 211.435 122.810 211.575 ;
        RECT 105.545 211.295 105.835 211.390 ;
        RECT 95.825 211.095 97.880 211.235 ;
        RECT 99.050 211.235 99.340 211.280 ;
        RECT 100.885 211.235 101.175 211.280 ;
        RECT 104.465 211.235 104.755 211.280 ;
        RECT 99.050 211.095 104.755 211.235 ;
        RECT 95.825 211.050 96.115 211.095 ;
        RECT 99.050 211.050 99.340 211.095 ;
        RECT 100.885 211.050 101.175 211.095 ;
        RECT 104.465 211.050 104.755 211.095 ;
        RECT 105.470 211.075 105.835 211.295 ;
        RECT 107.785 211.235 108.075 211.280 ;
        RECT 108.230 211.235 108.550 211.295 ;
        RECT 107.785 211.095 108.550 211.235 ;
        RECT 105.470 211.035 105.790 211.075 ;
        RECT 107.785 211.050 108.075 211.095 ;
        RECT 108.230 211.035 108.550 211.095 ;
        RECT 118.350 211.035 118.670 211.295 ;
        RECT 120.190 211.235 120.510 211.295 ;
        RECT 120.740 211.235 120.880 211.435 ;
        RECT 122.490 211.375 122.810 211.435 ;
        RECT 120.190 211.095 120.880 211.235 ;
        RECT 120.190 211.035 120.510 211.095 ;
        RECT 121.110 211.035 121.430 211.295 ;
        RECT 123.500 211.280 123.640 211.775 ;
        RECT 124.790 211.715 125.110 211.775 ;
        RECT 132.610 211.715 132.930 211.775 ;
        RECT 133.070 211.715 133.390 211.975 ;
        RECT 135.385 211.915 135.675 211.960 ;
        RECT 138.590 211.915 138.910 211.975 ;
        RECT 135.385 211.775 138.910 211.915 ;
        RECT 135.385 211.730 135.675 211.775 ;
        RECT 138.590 211.715 138.910 211.775 ;
        RECT 145.490 211.715 145.810 211.975 ;
        RECT 125.250 211.375 125.570 211.635 ;
        RECT 127.545 211.575 128.195 211.620 ;
        RECT 128.930 211.575 129.250 211.635 ;
        RECT 131.145 211.575 131.435 211.620 ;
        RECT 127.545 211.435 131.435 211.575 ;
        RECT 127.545 211.390 128.195 211.435 ;
        RECT 128.930 211.375 129.250 211.435 ;
        RECT 130.845 211.390 131.435 211.435 ;
        RECT 134.925 211.575 135.215 211.620 ;
        RECT 139.970 211.575 140.290 211.635 ;
        RECT 134.925 211.435 140.290 211.575 ;
        RECT 134.925 211.390 135.215 211.435 ;
        RECT 123.425 211.050 123.715 211.280 ;
        RECT 124.350 211.235 124.640 211.280 ;
        RECT 126.185 211.235 126.475 211.280 ;
        RECT 129.765 211.235 130.055 211.280 ;
        RECT 124.350 211.095 130.055 211.235 ;
        RECT 124.350 211.050 124.640 211.095 ;
        RECT 126.185 211.050 126.475 211.095 ;
        RECT 129.765 211.050 130.055 211.095 ;
        RECT 130.845 211.075 131.135 211.390 ;
        RECT 72.900 210.755 76.260 210.895 ;
        RECT 39.690 210.555 40.010 210.615 ;
        RECT 55.330 210.555 55.650 210.615 ;
        RECT 59.485 210.555 59.775 210.600 ;
        RECT 71.890 210.555 72.210 210.615 ;
        RECT 31.870 210.415 40.010 210.555 ;
        RECT 26.350 210.355 26.670 210.415 ;
        RECT 31.870 210.355 32.190 210.415 ;
        RECT 39.690 210.355 40.010 210.415 ;
        RECT 45.760 210.415 55.105 210.555 ;
        RECT 39.230 210.215 39.550 210.275 ;
        RECT 45.760 210.215 45.900 210.415 ;
        RECT 39.230 210.075 45.900 210.215 ;
        RECT 46.605 210.215 46.895 210.260 ;
        RECT 47.510 210.215 47.830 210.275 ;
        RECT 46.605 210.075 47.830 210.215 ;
        RECT 39.230 210.015 39.550 210.075 ;
        RECT 46.605 210.030 46.895 210.075 ;
        RECT 47.510 210.015 47.830 210.075 ;
        RECT 51.190 210.215 51.510 210.275 ;
        RECT 51.665 210.215 51.955 210.260 ;
        RECT 51.190 210.075 51.955 210.215 ;
        RECT 51.190 210.015 51.510 210.075 ;
        RECT 51.665 210.030 51.955 210.075 ;
        RECT 53.030 210.215 53.350 210.275 ;
        RECT 53.505 210.215 53.795 210.260 ;
        RECT 53.030 210.075 53.795 210.215 ;
        RECT 54.965 210.215 55.105 210.415 ;
        RECT 55.330 210.415 72.210 210.555 ;
        RECT 72.440 210.555 72.580 210.710 ;
        RECT 78.330 210.695 78.650 210.955 ;
        RECT 78.790 210.695 79.110 210.955 ;
        RECT 86.150 210.695 86.470 210.955 ;
        RECT 88.450 210.895 88.770 210.955 ;
        RECT 98.585 210.895 98.875 210.940 ;
        RECT 105.560 210.895 105.700 211.035 ;
        RECT 88.450 210.755 98.875 210.895 ;
        RECT 88.450 210.695 88.770 210.755 ;
        RECT 80.170 210.555 80.490 210.615 ;
        RECT 72.440 210.415 80.490 210.555 ;
        RECT 55.330 210.355 55.650 210.415 ;
        RECT 59.485 210.370 59.775 210.415 ;
        RECT 71.890 210.355 72.210 210.415 ;
        RECT 80.170 210.355 80.490 210.415 ;
        RECT 81.090 210.555 81.410 210.615 ;
        RECT 88.910 210.555 89.230 210.615 ;
        RECT 81.090 210.415 89.230 210.555 ;
        RECT 81.090 210.355 81.410 210.415 ;
        RECT 88.910 210.355 89.230 210.415 ;
        RECT 89.845 210.555 90.135 210.600 ;
        RECT 91.685 210.555 91.975 210.600 ;
        RECT 89.845 210.415 91.975 210.555 ;
        RECT 89.845 210.370 90.135 210.415 ;
        RECT 91.685 210.370 91.975 210.415 ;
        RECT 69.130 210.215 69.450 210.275 ;
        RECT 54.965 210.075 69.450 210.215 ;
        RECT 53.030 210.015 53.350 210.075 ;
        RECT 53.505 210.030 53.795 210.075 ;
        RECT 69.130 210.015 69.450 210.075 ;
        RECT 70.050 210.215 70.370 210.275 ;
        RECT 73.745 210.215 74.035 210.260 ;
        RECT 70.050 210.075 74.035 210.215 ;
        RECT 70.050 210.015 70.370 210.075 ;
        RECT 73.745 210.030 74.035 210.075 ;
        RECT 76.030 210.015 76.350 210.275 ;
        RECT 82.010 210.215 82.330 210.275 ;
        RECT 82.485 210.215 82.775 210.260 ;
        RECT 82.010 210.075 82.775 210.215 ;
        RECT 82.010 210.015 82.330 210.075 ;
        RECT 82.485 210.030 82.775 210.075 ;
        RECT 82.930 210.215 83.250 210.275 ;
        RECT 83.865 210.215 84.155 210.260 ;
        RECT 82.930 210.075 84.155 210.215 ;
        RECT 82.930 210.015 83.250 210.075 ;
        RECT 83.865 210.030 84.155 210.075 ;
        RECT 84.770 210.215 85.090 210.275 ;
        RECT 86.610 210.215 86.930 210.275 ;
        RECT 84.770 210.075 86.930 210.215 ;
        RECT 84.770 210.015 85.090 210.075 ;
        RECT 86.610 210.015 86.930 210.075 ;
        RECT 90.750 210.215 91.070 210.275 ;
        RECT 93.970 210.215 94.290 210.275 ;
        RECT 96.745 210.215 97.035 210.260 ;
        RECT 90.750 210.075 97.035 210.215 ;
        RECT 97.740 210.215 97.880 210.755 ;
        RECT 98.585 210.710 98.875 210.755 ;
        RECT 99.120 210.755 105.700 210.895 ;
        RECT 98.110 210.555 98.430 210.615 ;
        RECT 99.120 210.555 99.260 210.755 ;
        RECT 116.525 210.710 116.815 210.940 ;
        RECT 117.430 210.895 117.750 210.955 ;
        RECT 119.745 210.895 120.035 210.940 ;
        RECT 117.430 210.755 120.035 210.895 ;
        RECT 98.110 210.415 99.260 210.555 ;
        RECT 99.455 210.555 99.745 210.600 ;
        RECT 101.345 210.555 101.635 210.600 ;
        RECT 104.465 210.555 104.755 210.600 ;
        RECT 99.455 210.415 104.755 210.555 ;
        RECT 98.110 210.355 98.430 210.415 ;
        RECT 99.455 210.370 99.745 210.415 ;
        RECT 101.345 210.370 101.635 210.415 ;
        RECT 104.465 210.370 104.755 210.415 ;
        RECT 107.770 210.555 108.090 210.615 ;
        RECT 116.600 210.555 116.740 210.710 ;
        RECT 117.430 210.695 117.750 210.755 ;
        RECT 119.745 210.710 120.035 210.755 ;
        RECT 120.650 210.695 120.970 210.955 ;
        RECT 123.885 210.710 124.175 210.940 ;
        RECT 127.550 210.895 127.870 210.955 ;
        RECT 135.000 210.895 135.140 211.390 ;
        RECT 139.970 211.375 140.290 211.435 ;
        RECT 135.370 211.235 135.690 211.295 ;
        RECT 140.905 211.235 141.195 211.280 ;
        RECT 135.370 211.095 141.195 211.235 ;
        RECT 135.370 211.035 135.690 211.095 ;
        RECT 140.905 211.050 141.195 211.095 ;
        RECT 144.570 211.035 144.890 211.295 ;
        RECT 127.550 210.755 135.140 210.895 ;
        RECT 135.830 210.895 136.150 210.955 ;
        RECT 139.970 210.895 140.290 210.955 ;
        RECT 135.830 210.755 140.290 210.895 ;
        RECT 123.960 210.555 124.100 210.710 ;
        RECT 127.550 210.695 127.870 210.755 ;
        RECT 135.830 210.695 136.150 210.755 ;
        RECT 139.970 210.695 140.290 210.755 ;
        RECT 107.770 210.415 124.100 210.555 ;
        RECT 107.770 210.355 108.090 210.415 ;
        RECT 107.860 210.215 108.000 210.355 ;
        RECT 97.740 210.075 108.000 210.215 ;
        RECT 117.905 210.215 118.195 210.260 ;
        RECT 119.270 210.215 119.590 210.275 ;
        RECT 117.905 210.075 119.590 210.215 ;
        RECT 90.750 210.015 91.070 210.075 ;
        RECT 93.970 210.015 94.290 210.075 ;
        RECT 96.745 210.030 97.035 210.075 ;
        RECT 117.905 210.030 118.195 210.075 ;
        RECT 119.270 210.015 119.590 210.075 ;
        RECT 119.730 210.215 120.050 210.275 ;
        RECT 122.965 210.215 123.255 210.260 ;
        RECT 119.730 210.075 123.255 210.215 ;
        RECT 123.960 210.215 124.100 210.415 ;
        RECT 124.755 210.555 125.045 210.600 ;
        RECT 126.645 210.555 126.935 210.600 ;
        RECT 129.765 210.555 130.055 210.600 ;
        RECT 124.755 210.415 130.055 210.555 ;
        RECT 124.755 210.370 125.045 210.415 ;
        RECT 126.645 210.370 126.935 210.415 ;
        RECT 129.765 210.370 130.055 210.415 ;
        RECT 130.310 210.215 130.630 210.275 ;
        RECT 123.960 210.075 130.630 210.215 ;
        RECT 119.730 210.015 120.050 210.075 ;
        RECT 122.965 210.030 123.255 210.075 ;
        RECT 130.310 210.015 130.630 210.075 ;
        RECT 132.625 210.215 132.915 210.260 ;
        RECT 134.450 210.215 134.770 210.275 ;
        RECT 132.625 210.075 134.770 210.215 ;
        RECT 132.625 210.030 132.915 210.075 ;
        RECT 134.450 210.015 134.770 210.075 ;
        RECT 141.810 210.015 142.130 210.275 ;
        RECT 13.860 209.395 147.720 209.875 ;
        RECT 27.270 208.995 27.590 209.255 ;
        RECT 30.490 209.195 30.810 209.255 ;
        RECT 35.090 209.195 35.410 209.255 ;
        RECT 30.490 209.055 35.410 209.195 ;
        RECT 30.490 208.995 30.810 209.055 ;
        RECT 35.090 208.995 35.410 209.055 ;
        RECT 35.550 209.195 35.870 209.255 ;
        RECT 36.945 209.195 37.235 209.240 ;
        RECT 35.550 209.055 37.235 209.195 ;
        RECT 35.550 208.995 35.870 209.055 ;
        RECT 36.945 209.010 37.235 209.055 ;
        RECT 37.390 209.195 37.710 209.255 ;
        RECT 37.390 209.055 38.540 209.195 ;
        RECT 37.390 208.995 37.710 209.055 ;
        RECT 14.170 208.855 14.490 208.915 ;
        RECT 15.785 208.855 16.075 208.900 ;
        RECT 14.170 208.715 16.075 208.855 ;
        RECT 14.170 208.655 14.490 208.715 ;
        RECT 15.785 208.670 16.075 208.715 ;
        RECT 24.065 208.855 24.355 208.900 ;
        RECT 27.730 208.855 28.050 208.915 ;
        RECT 33.250 208.855 33.570 208.915 ;
        RECT 37.850 208.855 38.170 208.915 ;
        RECT 24.065 208.715 28.050 208.855 ;
        RECT 24.065 208.670 24.355 208.715 ;
        RECT 27.730 208.655 28.050 208.715 ;
        RECT 29.200 208.715 33.570 208.855 ;
        RECT 28.650 208.515 28.970 208.575 ;
        RECT 25.060 208.375 28.970 208.515 ;
        RECT 16.690 207.975 17.010 208.235 ;
        RECT 18.545 208.175 18.835 208.220 ;
        RECT 22.670 208.175 22.990 208.235 ;
        RECT 18.545 208.035 22.990 208.175 ;
        RECT 18.545 207.990 18.835 208.035 ;
        RECT 22.670 207.975 22.990 208.035 ;
        RECT 24.510 208.175 24.830 208.235 ;
        RECT 25.060 208.220 25.200 208.375 ;
        RECT 28.650 208.315 28.970 208.375 ;
        RECT 24.985 208.175 25.275 208.220 ;
        RECT 24.510 208.035 25.275 208.175 ;
        RECT 24.510 207.975 24.830 208.035 ;
        RECT 24.985 207.990 25.275 208.035 ;
        RECT 25.445 207.990 25.735 208.220 ;
        RECT 25.905 208.175 26.195 208.220 ;
        RECT 28.190 208.175 28.510 208.235 ;
        RECT 29.200 208.220 29.340 208.715 ;
        RECT 33.250 208.655 33.570 208.715 ;
        RECT 33.800 208.715 38.170 208.855 ;
        RECT 38.400 208.855 38.540 209.055 ;
        RECT 38.770 208.995 39.090 209.255 ;
        RECT 44.305 209.195 44.595 209.240 ;
        RECT 47.050 209.195 47.370 209.255 ;
        RECT 47.985 209.195 48.275 209.240 ;
        RECT 44.305 209.055 47.370 209.195 ;
        RECT 44.305 209.010 44.595 209.055 ;
        RECT 47.050 208.995 47.370 209.055 ;
        RECT 47.600 209.055 48.275 209.195 ;
        RECT 42.910 208.855 43.230 208.915 ;
        RECT 44.750 208.855 45.070 208.915 ;
        RECT 38.400 208.715 45.070 208.855 ;
        RECT 33.800 208.560 33.940 208.715 ;
        RECT 37.850 208.655 38.170 208.715 ;
        RECT 42.910 208.655 43.230 208.715 ;
        RECT 44.750 208.655 45.070 208.715 ;
        RECT 30.505 208.515 30.795 208.560 ;
        RECT 31.425 208.515 31.715 208.560 ;
        RECT 32.805 208.515 33.095 208.560 ;
        RECT 30.505 208.375 31.715 208.515 ;
        RECT 30.505 208.330 30.795 208.375 ;
        RECT 31.425 208.330 31.715 208.375 ;
        RECT 31.960 208.375 33.095 208.515 ;
        RECT 25.905 208.035 28.510 208.175 ;
        RECT 25.905 207.990 26.195 208.035 ;
        RECT 17.610 207.295 17.930 207.555 ;
        RECT 25.520 207.495 25.660 207.990 ;
        RECT 28.190 207.975 28.510 208.035 ;
        RECT 29.125 207.990 29.415 208.220 ;
        RECT 30.950 208.175 31.270 208.235 ;
        RECT 31.960 208.175 32.100 208.375 ;
        RECT 32.805 208.330 33.095 208.375 ;
        RECT 33.725 208.330 34.015 208.560 ;
        RECT 41.545 208.515 41.835 208.560 ;
        RECT 41.990 208.515 42.310 208.575 ;
        RECT 47.600 208.515 47.740 209.055 ;
        RECT 47.985 209.010 48.275 209.055 ;
        RECT 52.110 209.195 52.430 209.255 ;
        RECT 53.045 209.195 53.335 209.240 ;
        RECT 52.110 209.055 53.335 209.195 ;
        RECT 52.110 208.995 52.430 209.055 ;
        RECT 53.045 209.010 53.335 209.055 ;
        RECT 53.490 209.195 53.810 209.255 ;
        RECT 54.885 209.195 55.175 209.240 ;
        RECT 53.490 209.055 55.175 209.195 ;
        RECT 53.490 208.995 53.810 209.055 ;
        RECT 54.885 209.010 55.175 209.055 ;
        RECT 55.790 208.995 56.110 209.255 ;
        RECT 56.250 209.195 56.570 209.255 ;
        RECT 68.670 209.195 68.990 209.255 ;
        RECT 56.250 209.055 68.990 209.195 ;
        RECT 56.250 208.995 56.570 209.055 ;
        RECT 68.670 208.995 68.990 209.055 ;
        RECT 70.985 209.195 71.275 209.240 ;
        RECT 71.430 209.195 71.750 209.255 ;
        RECT 70.985 209.055 71.750 209.195 ;
        RECT 70.985 209.010 71.275 209.055 ;
        RECT 71.430 208.995 71.750 209.055 ;
        RECT 71.890 209.195 72.210 209.255 ;
        RECT 75.570 209.195 75.890 209.255 ;
        RECT 71.890 209.055 75.890 209.195 ;
        RECT 71.890 208.995 72.210 209.055 ;
        RECT 75.570 208.995 75.890 209.055 ;
        RECT 76.505 209.195 76.795 209.240 ;
        RECT 77.410 209.195 77.730 209.255 ;
        RECT 76.505 209.055 77.730 209.195 ;
        RECT 76.505 209.010 76.795 209.055 ;
        RECT 77.410 208.995 77.730 209.055 ;
        RECT 78.330 209.195 78.650 209.255 ;
        RECT 79.725 209.195 80.015 209.240 ;
        RECT 78.330 209.055 80.015 209.195 ;
        RECT 78.330 208.995 78.650 209.055 ;
        RECT 79.725 209.010 80.015 209.055 ;
        RECT 86.150 209.195 86.470 209.255 ;
        RECT 87.085 209.195 87.375 209.240 ;
        RECT 86.150 209.055 87.375 209.195 ;
        RECT 86.150 208.995 86.470 209.055 ;
        RECT 87.085 209.010 87.375 209.055 ;
        RECT 93.050 209.195 93.370 209.255 ;
        RECT 99.045 209.195 99.335 209.240 ;
        RECT 105.025 209.195 105.315 209.240 ;
        RECT 93.050 209.055 99.335 209.195 ;
        RECT 93.050 208.995 93.370 209.055 ;
        RECT 99.045 209.010 99.335 209.055 ;
        RECT 100.500 209.055 105.315 209.195 ;
        RECT 59.010 208.855 59.330 208.915 ;
        RECT 61.310 208.855 61.630 208.915 ;
        RECT 57.720 208.715 61.630 208.855 ;
        RECT 53.030 208.515 53.350 208.575 ;
        RECT 57.720 208.560 57.860 208.715 ;
        RECT 59.010 208.655 59.330 208.715 ;
        RECT 61.310 208.655 61.630 208.715 ;
        RECT 62.345 208.855 62.635 208.900 ;
        RECT 65.465 208.855 65.755 208.900 ;
        RECT 67.355 208.855 67.645 208.900 ;
        RECT 73.730 208.855 74.050 208.915 ;
        RECT 62.345 208.715 67.645 208.855 ;
        RECT 62.345 208.670 62.635 208.715 ;
        RECT 65.465 208.670 65.755 208.715 ;
        RECT 67.355 208.670 67.645 208.715 ;
        RECT 72.900 208.715 74.050 208.855 ;
        RECT 53.505 208.515 53.795 208.560 ;
        RECT 35.640 208.375 42.310 208.515 ;
        RECT 35.640 208.235 35.780 208.375 ;
        RECT 38.400 208.235 38.540 208.375 ;
        RECT 41.545 208.330 41.835 208.375 ;
        RECT 41.990 208.315 42.310 208.375 ;
        RECT 42.540 208.375 47.740 208.515 ;
        RECT 48.060 208.375 53.795 208.515 ;
        RECT 30.950 208.035 32.100 208.175 ;
        RECT 30.950 207.975 31.270 208.035 ;
        RECT 32.345 207.990 32.635 208.220 ;
        RECT 33.265 208.175 33.555 208.220 ;
        RECT 34.630 208.175 34.950 208.235 ;
        RECT 33.265 208.035 34.950 208.175 ;
        RECT 33.265 207.990 33.555 208.035 ;
        RECT 27.730 207.835 28.050 207.895 ;
        RECT 32.420 207.835 32.560 207.990 ;
        RECT 34.630 207.975 34.950 208.035 ;
        RECT 35.090 207.975 35.410 208.235 ;
        RECT 35.550 207.975 35.870 208.235 ;
        RECT 36.025 208.175 36.315 208.220 ;
        RECT 36.930 208.175 37.250 208.235 ;
        RECT 36.025 208.035 37.250 208.175 ;
        RECT 36.025 207.990 36.315 208.035 ;
        RECT 36.930 207.975 37.250 208.035 ;
        RECT 37.390 207.975 37.710 208.235 ;
        RECT 38.310 207.975 38.630 208.235 ;
        RECT 42.540 208.175 42.680 208.375 ;
        RECT 48.060 208.235 48.200 208.375 ;
        RECT 53.030 208.315 53.350 208.375 ;
        RECT 53.505 208.330 53.795 208.375 ;
        RECT 53.965 208.330 54.255 208.560 ;
        RECT 57.645 208.330 57.935 208.560 ;
        RECT 63.150 208.515 63.470 208.575 ;
        RECT 60.940 208.375 63.470 208.515 ;
        RECT 38.860 208.035 42.680 208.175 ;
        RECT 42.925 208.175 43.215 208.220 ;
        RECT 44.290 208.175 44.610 208.235 ;
        RECT 42.925 208.035 44.610 208.175 ;
        RECT 27.730 207.695 32.560 207.835 ;
        RECT 37.020 207.835 37.160 207.975 ;
        RECT 38.860 207.835 39.000 208.035 ;
        RECT 42.925 207.990 43.215 208.035 ;
        RECT 44.290 207.975 44.610 208.035 ;
        RECT 45.210 207.975 45.530 208.235 ;
        RECT 46.590 207.975 46.910 208.235 ;
        RECT 47.970 207.975 48.290 208.235 ;
        RECT 49.350 208.175 49.670 208.235 ;
        RECT 49.825 208.175 50.115 208.220 ;
        RECT 49.350 208.035 50.115 208.175 ;
        RECT 49.350 207.975 49.670 208.035 ;
        RECT 49.825 207.990 50.115 208.035 ;
        RECT 50.270 207.975 50.590 208.235 ;
        RECT 54.040 208.175 54.180 208.330 ;
        RECT 50.820 208.035 54.180 208.175 ;
        RECT 37.020 207.695 39.000 207.835 ;
        RECT 39.230 207.835 39.550 207.895 ;
        RECT 41.085 207.835 41.375 207.880 ;
        RECT 39.230 207.695 41.375 207.835 ;
        RECT 27.730 207.635 28.050 207.695 ;
        RECT 39.230 207.635 39.550 207.695 ;
        RECT 41.085 207.650 41.375 207.695 ;
        RECT 43.385 207.835 43.675 207.880 ;
        RECT 50.360 207.835 50.500 207.975 ;
        RECT 43.385 207.695 50.500 207.835 ;
        RECT 43.385 207.650 43.675 207.695 ;
        RECT 28.650 207.495 28.970 207.555 ;
        RECT 25.520 207.355 28.970 207.495 ;
        RECT 28.650 207.295 28.970 207.355 ;
        RECT 29.585 207.495 29.875 207.540 ;
        RECT 32.330 207.495 32.650 207.555 ;
        RECT 37.390 207.495 37.710 207.555 ;
        RECT 29.585 207.355 37.710 207.495 ;
        RECT 29.585 207.310 29.875 207.355 ;
        RECT 32.330 207.295 32.650 207.355 ;
        RECT 37.390 207.295 37.710 207.355 ;
        RECT 38.325 207.495 38.615 207.540 ;
        RECT 40.150 207.495 40.470 207.555 ;
        RECT 38.325 207.355 40.470 207.495 ;
        RECT 38.325 207.310 38.615 207.355 ;
        RECT 40.150 207.295 40.470 207.355 ;
        RECT 40.625 207.495 40.915 207.540 ;
        RECT 41.530 207.495 41.850 207.555 ;
        RECT 40.625 207.355 41.850 207.495 ;
        RECT 40.625 207.310 40.915 207.355 ;
        RECT 41.530 207.295 41.850 207.355 ;
        RECT 46.145 207.495 46.435 207.540 ;
        RECT 47.065 207.495 47.355 207.540 ;
        RECT 46.145 207.355 47.355 207.495 ;
        RECT 46.145 207.310 46.435 207.355 ;
        RECT 47.065 207.310 47.355 207.355 ;
        RECT 47.510 207.495 47.830 207.555 ;
        RECT 50.820 207.495 50.960 208.035 ;
        RECT 55.330 207.975 55.650 208.235 ;
        RECT 56.710 208.175 57.030 208.235 ;
        RECT 60.940 208.175 61.080 208.375 ;
        RECT 63.150 208.315 63.470 208.375 ;
        RECT 66.830 208.515 67.150 208.575 ;
        RECT 68.225 208.515 68.515 208.560 ;
        RECT 66.830 208.375 68.515 208.515 ;
        RECT 66.830 208.315 67.150 208.375 ;
        RECT 68.225 208.330 68.515 208.375 ;
        RECT 70.050 208.315 70.370 208.575 ;
        RECT 70.525 208.515 70.815 208.560 ;
        RECT 71.445 208.515 71.735 208.560 ;
        RECT 72.350 208.515 72.670 208.575 ;
        RECT 70.525 208.375 71.200 208.515 ;
        RECT 70.525 208.330 70.815 208.375 ;
        RECT 56.710 208.035 61.080 208.175 ;
        RECT 56.710 207.975 57.030 208.035 ;
        RECT 61.265 207.880 61.555 208.195 ;
        RECT 62.345 208.175 62.635 208.220 ;
        RECT 65.925 208.175 66.215 208.220 ;
        RECT 67.760 208.175 68.050 208.220 ;
        RECT 62.345 208.035 68.050 208.175 ;
        RECT 62.345 207.990 62.635 208.035 ;
        RECT 65.925 207.990 66.215 208.035 ;
        RECT 67.760 207.990 68.050 208.035 ;
        RECT 60.965 207.835 61.555 207.880 ;
        RECT 64.070 207.880 64.390 207.895 ;
        RECT 64.070 207.835 64.855 207.880 ;
        RECT 60.965 207.695 64.855 207.835 ;
        RECT 60.965 207.650 61.255 207.695 ;
        RECT 64.070 207.650 64.855 207.695 ;
        RECT 66.370 207.835 66.690 207.895 ;
        RECT 66.845 207.835 67.135 207.880 ;
        RECT 66.370 207.695 67.135 207.835 ;
        RECT 64.070 207.635 64.390 207.650 ;
        RECT 66.370 207.635 66.690 207.695 ;
        RECT 66.845 207.650 67.135 207.695 ;
        RECT 47.510 207.355 50.960 207.495 ;
        RECT 51.205 207.495 51.495 207.540 ;
        RECT 51.650 207.495 51.970 207.555 ;
        RECT 51.205 207.355 51.970 207.495 ;
        RECT 47.510 207.295 47.830 207.355 ;
        RECT 51.205 207.310 51.495 207.355 ;
        RECT 51.650 207.295 51.970 207.355 ;
        RECT 59.470 207.295 59.790 207.555 ;
        RECT 71.060 207.495 71.200 208.375 ;
        RECT 71.445 208.375 72.670 208.515 ;
        RECT 71.445 208.330 71.735 208.375 ;
        RECT 72.350 208.315 72.670 208.375 ;
        RECT 71.905 208.175 72.195 208.220 ;
        RECT 72.900 208.175 73.040 208.715 ;
        RECT 73.730 208.655 74.050 208.715 ;
        RECT 74.190 208.855 74.510 208.915 ;
        RECT 76.030 208.855 76.350 208.915 ;
        RECT 90.750 208.855 91.070 208.915 ;
        RECT 74.190 208.715 76.350 208.855 ;
        RECT 74.190 208.655 74.510 208.715 ;
        RECT 76.030 208.655 76.350 208.715 ;
        RECT 84.860 208.715 91.070 208.855 ;
        RECT 73.285 208.515 73.575 208.560 ;
        RECT 73.285 208.375 76.720 208.515 ;
        RECT 73.285 208.330 73.575 208.375 ;
        RECT 71.905 208.035 73.040 208.175 ;
        RECT 71.905 207.990 72.195 208.035 ;
        RECT 73.745 207.990 74.035 208.220 ;
        RECT 74.205 207.990 74.495 208.220 ;
        RECT 74.665 208.175 74.955 208.220 ;
        RECT 75.110 208.175 75.430 208.235 ;
        RECT 74.665 208.035 75.430 208.175 ;
        RECT 74.665 207.990 74.955 208.035 ;
        RECT 72.365 207.495 72.655 207.540 ;
        RECT 71.060 207.355 72.655 207.495 ;
        RECT 72.365 207.310 72.655 207.355 ;
        RECT 73.270 207.495 73.590 207.555 ;
        RECT 73.820 207.495 73.960 207.990 ;
        RECT 74.280 207.555 74.420 207.990 ;
        RECT 75.110 207.975 75.430 208.035 ;
        RECT 75.570 207.975 75.890 208.235 ;
        RECT 76.580 208.175 76.720 208.375 ;
        RECT 76.950 208.315 77.270 208.575 ;
        RECT 82.930 208.315 83.250 208.575 ;
        RECT 84.860 208.560 85.000 208.715 ;
        RECT 90.750 208.655 91.070 208.715 ;
        RECT 95.365 208.670 95.655 208.900 ;
        RECT 95.810 208.855 96.130 208.915 ;
        RECT 98.570 208.855 98.890 208.915 ;
        RECT 100.500 208.855 100.640 209.055 ;
        RECT 105.025 209.010 105.315 209.055 ;
        RECT 106.850 209.195 107.170 209.255 ;
        RECT 107.325 209.195 107.615 209.240 ;
        RECT 125.710 209.195 126.030 209.255 ;
        RECT 129.850 209.195 130.170 209.255 ;
        RECT 106.850 209.055 107.615 209.195 ;
        RECT 106.850 208.995 107.170 209.055 ;
        RECT 107.325 209.010 107.615 209.055 ;
        RECT 108.320 209.055 130.170 209.195 ;
        RECT 95.810 208.715 98.890 208.855 ;
        RECT 84.785 208.330 85.075 208.560 ;
        RECT 85.690 208.515 86.010 208.575 ;
        RECT 86.165 208.515 86.455 208.560 ;
        RECT 85.690 208.375 86.455 208.515 ;
        RECT 85.690 208.315 86.010 208.375 ;
        RECT 86.165 208.330 86.455 208.375 ;
        RECT 87.070 208.515 87.390 208.575 ;
        RECT 95.440 208.515 95.580 208.670 ;
        RECT 95.810 208.655 96.130 208.715 ;
        RECT 98.570 208.655 98.890 208.715 ;
        RECT 99.120 208.715 100.640 208.855 ;
        RECT 99.120 208.515 99.260 208.715 ;
        RECT 87.070 208.375 89.140 208.515 ;
        RECT 87.070 208.315 87.390 208.375 ;
        RECT 78.790 208.175 79.110 208.235 ;
        RECT 76.580 208.035 79.110 208.175 ;
        RECT 78.790 207.975 79.110 208.035 ;
        RECT 80.630 207.975 80.950 208.235 ;
        RECT 81.090 207.975 81.410 208.235 ;
        RECT 83.850 208.175 84.170 208.235 ;
        RECT 85.245 208.175 85.535 208.220 ;
        RECT 83.850 208.035 85.535 208.175 ;
        RECT 83.850 207.975 84.170 208.035 ;
        RECT 85.245 207.990 85.535 208.035 ;
        RECT 86.625 208.175 86.915 208.220 ;
        RECT 87.530 208.175 87.850 208.235 ;
        RECT 86.625 208.035 87.850 208.175 ;
        RECT 86.625 207.990 86.915 208.035 ;
        RECT 87.530 207.975 87.850 208.035 ;
        RECT 87.990 207.975 88.310 208.235 ;
        RECT 88.450 207.975 88.770 208.235 ;
        RECT 89.000 208.220 89.140 208.375 ;
        RECT 89.590 208.375 91.900 208.515 ;
        RECT 89.590 208.220 89.730 208.375 ;
        RECT 88.925 207.990 89.215 208.220 ;
        RECT 89.515 207.990 89.805 208.220 ;
        RECT 90.305 208.175 90.595 208.220 ;
        RECT 91.210 208.175 91.530 208.235 ;
        RECT 90.305 208.035 91.530 208.175 ;
        RECT 91.760 208.175 91.900 208.375 ;
        RECT 93.140 208.375 95.580 208.515 ;
        RECT 96.820 208.375 99.260 208.515 ;
        RECT 93.140 208.175 93.280 208.375 ;
        RECT 91.760 208.035 93.280 208.175 ;
        RECT 90.305 207.990 90.595 208.035 ;
        RECT 91.210 207.975 91.530 208.035 ;
        RECT 94.890 207.975 95.210 208.235 ;
        RECT 96.820 208.175 96.960 208.375 ;
        RECT 99.950 208.315 100.270 208.575 ;
        RECT 100.500 208.560 100.640 208.715 ;
        RECT 100.870 208.855 101.190 208.915 ;
        RECT 108.320 208.855 108.460 209.055 ;
        RECT 125.710 208.995 126.030 209.055 ;
        RECT 129.850 208.995 130.170 209.055 ;
        RECT 145.490 208.995 145.810 209.255 ;
        RECT 100.870 208.715 108.460 208.855 ;
        RECT 108.655 208.855 108.945 208.900 ;
        RECT 110.545 208.855 110.835 208.900 ;
        RECT 113.665 208.855 113.955 208.900 ;
        RECT 108.655 208.715 113.955 208.855 ;
        RECT 100.870 208.655 101.190 208.715 ;
        RECT 100.425 208.330 100.715 208.560 ;
        RECT 95.440 208.035 96.960 208.175 ;
        RECT 97.205 208.175 97.495 208.220 ;
        RECT 97.650 208.175 97.970 208.235 ;
        RECT 97.205 208.035 97.970 208.175 ;
        RECT 78.330 207.835 78.650 207.895 ;
        RECT 79.710 207.835 80.030 207.895 ;
        RECT 78.330 207.695 80.030 207.835 ;
        RECT 78.330 207.635 78.650 207.695 ;
        RECT 79.710 207.635 80.030 207.695 ;
        RECT 81.550 207.635 81.870 207.895 ;
        RECT 92.590 207.880 92.910 207.895 ;
        RECT 82.255 207.835 82.545 207.880 ;
        RECT 82.255 207.695 87.300 207.835 ;
        RECT 82.255 207.650 82.545 207.695 ;
        RECT 73.270 207.355 73.960 207.495 ;
        RECT 74.190 207.495 74.510 207.555 ;
        RECT 79.250 207.495 79.570 207.555 ;
        RECT 74.190 207.355 79.570 207.495 ;
        RECT 73.270 207.295 73.590 207.355 ;
        RECT 74.190 207.295 74.510 207.355 ;
        RECT 79.250 207.295 79.570 207.355 ;
        RECT 84.785 207.495 85.075 207.540 ;
        RECT 86.150 207.495 86.470 207.555 ;
        RECT 84.785 207.355 86.470 207.495 ;
        RECT 87.160 207.495 87.300 207.695 ;
        RECT 92.480 207.650 92.910 207.880 ;
        RECT 93.065 207.835 93.355 207.880 ;
        RECT 93.970 207.835 94.290 207.895 ;
        RECT 93.065 207.695 94.290 207.835 ;
        RECT 93.065 207.650 93.355 207.695 ;
        RECT 92.590 207.635 92.910 207.650 ;
        RECT 93.970 207.635 94.290 207.695 ;
        RECT 94.430 207.835 94.750 207.895 ;
        RECT 95.440 207.835 95.580 208.035 ;
        RECT 97.205 207.990 97.495 208.035 ;
        RECT 97.650 207.975 97.970 208.035 ;
        RECT 98.585 208.175 98.875 208.220 ;
        RECT 99.030 208.175 99.350 208.235 ;
        RECT 98.585 208.035 99.350 208.175 ;
        RECT 98.585 207.990 98.875 208.035 ;
        RECT 99.030 207.975 99.350 208.035 ;
        RECT 99.490 208.175 99.810 208.235 ;
        RECT 100.885 208.175 101.175 208.220 ;
        RECT 99.490 208.035 101.175 208.175 ;
        RECT 99.490 207.975 99.810 208.035 ;
        RECT 100.885 207.990 101.175 208.035 ;
        RECT 101.345 208.175 101.635 208.220 ;
        RECT 102.250 208.175 102.570 208.235 ;
        RECT 102.800 208.220 102.940 208.715 ;
        RECT 108.655 208.670 108.945 208.715 ;
        RECT 110.545 208.670 110.835 208.715 ;
        RECT 113.665 208.670 113.955 208.715 ;
        RECT 121.535 208.855 121.825 208.900 ;
        RECT 123.425 208.855 123.715 208.900 ;
        RECT 126.545 208.855 126.835 208.900 ;
        RECT 121.535 208.715 126.835 208.855 ;
        RECT 121.535 208.670 121.825 208.715 ;
        RECT 123.425 208.670 123.715 208.715 ;
        RECT 126.545 208.670 126.835 208.715 ;
        RECT 127.090 208.855 127.410 208.915 ;
        RECT 129.390 208.855 129.710 208.915 ;
        RECT 131.195 208.855 131.485 208.900 ;
        RECT 133.085 208.855 133.375 208.900 ;
        RECT 136.205 208.855 136.495 208.900 ;
        RECT 127.090 208.715 131.000 208.855 ;
        RECT 127.090 208.655 127.410 208.715 ;
        RECT 129.390 208.655 129.710 208.715 ;
        RECT 104.090 208.515 104.410 208.575 ;
        RECT 105.945 208.515 106.235 208.560 ;
        RECT 120.665 208.515 120.955 208.560 ;
        RECT 130.310 208.515 130.630 208.575 ;
        RECT 104.090 208.375 106.235 208.515 ;
        RECT 104.090 208.315 104.410 208.375 ;
        RECT 105.945 208.330 106.235 208.375 ;
        RECT 106.480 208.375 118.120 208.515 ;
        RECT 101.345 208.035 102.570 208.175 ;
        RECT 101.345 207.990 101.635 208.035 ;
        RECT 102.250 207.975 102.570 208.035 ;
        RECT 102.725 207.990 103.015 208.220 ;
        RECT 104.565 208.175 104.855 208.220 ;
        RECT 105.010 208.175 105.330 208.235 ;
        RECT 104.565 208.035 105.330 208.175 ;
        RECT 104.565 207.990 104.855 208.035 ;
        RECT 105.010 207.975 105.330 208.035 ;
        RECT 96.270 207.880 96.590 207.895 ;
        RECT 94.430 207.695 95.580 207.835 ;
        RECT 94.430 207.635 94.750 207.695 ;
        RECT 96.160 207.650 96.590 207.880 ;
        RECT 96.270 207.635 96.590 207.650 ;
        RECT 103.630 207.835 103.950 207.895 ;
        RECT 106.480 207.835 106.620 208.375 ;
        RECT 107.770 207.975 108.090 208.235 ;
        RECT 108.250 208.175 108.540 208.220 ;
        RECT 110.085 208.175 110.375 208.220 ;
        RECT 113.665 208.175 113.955 208.220 ;
        RECT 108.250 208.035 113.955 208.175 ;
        RECT 108.250 207.990 108.540 208.035 ;
        RECT 110.085 207.990 110.375 208.035 ;
        RECT 113.665 207.990 113.955 208.035 ;
        RECT 103.630 207.695 106.620 207.835 ;
        RECT 103.630 207.635 103.950 207.695 ;
        RECT 109.150 207.635 109.470 207.895 ;
        RECT 114.745 207.880 115.035 208.195 ;
        RECT 116.510 208.175 116.830 208.235 ;
        RECT 117.980 208.220 118.120 208.375 ;
        RECT 120.665 208.375 130.630 208.515 ;
        RECT 130.860 208.515 131.000 208.715 ;
        RECT 131.195 208.715 136.495 208.855 ;
        RECT 131.195 208.670 131.485 208.715 ;
        RECT 133.085 208.670 133.375 208.715 ;
        RECT 136.205 208.670 136.495 208.715 ;
        RECT 143.650 208.655 143.970 208.915 ;
        RECT 131.705 208.515 131.995 208.560 ;
        RECT 130.860 208.375 131.995 208.515 ;
        RECT 120.665 208.330 120.955 208.375 ;
        RECT 130.310 208.315 130.630 208.375 ;
        RECT 131.705 208.330 131.995 208.375 ;
        RECT 133.530 208.515 133.850 208.575 ;
        RECT 133.530 208.375 142.960 208.515 ;
        RECT 133.530 208.315 133.850 208.375 ;
        RECT 116.985 208.175 117.275 208.220 ;
        RECT 116.510 208.035 117.275 208.175 ;
        RECT 116.510 207.975 116.830 208.035 ;
        RECT 116.985 207.990 117.275 208.035 ;
        RECT 117.905 207.990 118.195 208.220 ;
        RECT 118.365 207.990 118.655 208.220 ;
        RECT 111.445 207.835 112.095 207.880 ;
        RECT 114.745 207.835 115.335 207.880 ;
        RECT 115.590 207.835 115.910 207.895 ;
        RECT 117.430 207.835 117.750 207.895 ;
        RECT 118.440 207.835 118.580 207.990 ;
        RECT 118.810 207.975 119.130 208.235 ;
        RECT 121.130 208.175 121.420 208.220 ;
        RECT 122.965 208.175 123.255 208.220 ;
        RECT 126.545 208.175 126.835 208.220 ;
        RECT 121.130 208.035 126.835 208.175 ;
        RECT 121.130 207.990 121.420 208.035 ;
        RECT 122.965 207.990 123.255 208.035 ;
        RECT 126.545 207.990 126.835 208.035 ;
        RECT 111.445 207.695 115.910 207.835 ;
        RECT 111.445 207.650 112.095 207.695 ;
        RECT 115.045 207.650 115.335 207.695 ;
        RECT 115.590 207.635 115.910 207.695 ;
        RECT 116.140 207.695 117.200 207.835 ;
        RECT 91.685 207.495 91.975 207.540 ;
        RECT 87.160 207.355 91.975 207.495 ;
        RECT 84.785 207.310 85.075 207.355 ;
        RECT 86.150 207.295 86.470 207.355 ;
        RECT 91.685 207.310 91.975 207.355 ;
        RECT 93.510 207.295 93.830 207.555 ;
        RECT 94.060 207.495 94.200 207.635 ;
        RECT 96.745 207.495 97.035 207.540 ;
        RECT 99.490 207.495 99.810 207.555 ;
        RECT 94.060 207.355 99.810 207.495 ;
        RECT 96.745 207.310 97.035 207.355 ;
        RECT 99.490 207.295 99.810 207.355 ;
        RECT 104.090 207.495 104.410 207.555 ;
        RECT 105.010 207.495 105.330 207.555 ;
        RECT 116.140 207.495 116.280 207.695 ;
        RECT 104.090 207.355 116.280 207.495 ;
        RECT 104.090 207.295 104.410 207.355 ;
        RECT 105.010 207.295 105.330 207.355 ;
        RECT 116.510 207.295 116.830 207.555 ;
        RECT 117.060 207.495 117.200 207.695 ;
        RECT 117.430 207.695 118.580 207.835 ;
        RECT 118.900 207.835 119.040 207.975 ;
        RECT 121.570 207.835 121.890 207.895 ;
        RECT 127.625 207.880 127.915 208.195 ;
        RECT 130.790 208.175 131.080 208.220 ;
        RECT 132.625 208.175 132.915 208.220 ;
        RECT 136.205 208.175 136.495 208.220 ;
        RECT 130.790 208.035 136.495 208.175 ;
        RECT 130.790 207.990 131.080 208.035 ;
        RECT 132.625 207.990 132.915 208.035 ;
        RECT 136.205 207.990 136.495 208.035 ;
        RECT 118.900 207.695 121.890 207.835 ;
        RECT 117.430 207.635 117.750 207.695 ;
        RECT 121.570 207.635 121.890 207.695 ;
        RECT 122.045 207.650 122.335 207.880 ;
        RECT 124.325 207.835 124.975 207.880 ;
        RECT 127.625 207.835 128.215 207.880 ;
        RECT 128.930 207.835 129.250 207.895 ;
        RECT 133.990 207.880 134.310 207.895 ;
        RECT 137.285 207.880 137.575 208.195 ;
        RECT 139.510 208.175 139.830 208.235 ;
        RECT 142.820 208.220 142.960 208.375 ;
        RECT 140.905 208.175 141.195 208.220 ;
        RECT 139.510 208.035 141.195 208.175 ;
        RECT 139.510 207.975 139.830 208.035 ;
        RECT 140.905 207.990 141.195 208.035 ;
        RECT 142.745 207.990 143.035 208.220 ;
        RECT 144.570 207.975 144.890 208.235 ;
        RECT 133.985 207.835 134.635 207.880 ;
        RECT 137.285 207.835 137.875 207.880 ;
        RECT 124.325 207.695 137.875 207.835 ;
        RECT 124.325 207.650 124.975 207.695 ;
        RECT 127.925 207.650 128.215 207.695 ;
        RECT 119.270 207.495 119.590 207.555 ;
        RECT 117.060 207.355 119.590 207.495 ;
        RECT 119.270 207.295 119.590 207.355 ;
        RECT 120.190 207.295 120.510 207.555 ;
        RECT 122.120 207.495 122.260 207.650 ;
        RECT 128.930 207.635 129.250 207.695 ;
        RECT 133.985 207.650 134.635 207.695 ;
        RECT 137.585 207.650 137.875 207.695 ;
        RECT 133.990 207.635 134.310 207.650 ;
        RECT 127.090 207.495 127.410 207.555 ;
        RECT 122.120 207.355 127.410 207.495 ;
        RECT 127.090 207.295 127.410 207.355 ;
        RECT 129.405 207.495 129.695 207.540 ;
        RECT 132.610 207.495 132.930 207.555 ;
        RECT 135.370 207.495 135.690 207.555 ;
        RECT 129.405 207.355 135.690 207.495 ;
        RECT 129.405 207.310 129.695 207.355 ;
        RECT 132.610 207.295 132.930 207.355 ;
        RECT 135.370 207.295 135.690 207.355 ;
        RECT 139.050 207.295 139.370 207.555 ;
        RECT 141.810 207.295 142.130 207.555 ;
        RECT 13.860 206.675 147.720 207.155 ;
        RECT 14.090 206.475 14.410 206.535 ;
        RECT 15.785 206.475 16.075 206.520 ;
        RECT 36.930 206.475 37.250 206.535 ;
        RECT 14.090 206.335 16.075 206.475 ;
        RECT 14.090 206.275 14.410 206.335 ;
        RECT 15.785 206.290 16.075 206.335 ;
        RECT 28.740 206.335 37.250 206.475 ;
        RECT 27.270 206.135 27.590 206.195 ;
        RECT 24.600 205.995 27.590 206.135 ;
        RECT 16.705 205.610 16.995 205.840 ;
        RECT 18.545 205.610 18.835 205.840 ;
        RECT 16.780 205.115 16.920 205.610 ;
        RECT 18.620 205.455 18.760 205.610 ;
        RECT 19.910 205.595 20.230 205.855 ;
        RECT 24.600 205.840 24.740 205.995 ;
        RECT 27.270 205.935 27.590 205.995 ;
        RECT 24.525 205.610 24.815 205.840 ;
        RECT 25.430 205.595 25.750 205.855 ;
        RECT 26.810 205.595 27.130 205.855 ;
        RECT 28.190 205.795 28.510 205.855 ;
        RECT 28.740 205.840 28.880 206.335 ;
        RECT 29.110 206.135 29.430 206.195 ;
        RECT 29.110 205.995 34.860 206.135 ;
        RECT 29.110 205.935 29.430 205.995 ;
        RECT 28.665 205.795 28.955 205.840 ;
        RECT 31.410 205.795 31.730 205.855 ;
        RECT 28.190 205.655 28.955 205.795 ;
        RECT 28.190 205.595 28.510 205.655 ;
        RECT 28.665 205.610 28.955 205.655 ;
        RECT 29.200 205.655 31.730 205.795 ;
        RECT 24.050 205.455 24.370 205.515 ;
        RECT 18.620 205.315 24.370 205.455 ;
        RECT 24.050 205.255 24.370 205.315 ;
        RECT 25.905 205.455 26.195 205.500 ;
        RECT 29.200 205.455 29.340 205.655 ;
        RECT 31.410 205.595 31.730 205.655 ;
        RECT 31.885 205.795 32.175 205.840 ;
        RECT 32.330 205.795 32.650 205.855 ;
        RECT 31.885 205.655 32.650 205.795 ;
        RECT 31.885 205.610 32.175 205.655 ;
        RECT 32.330 205.595 32.650 205.655 ;
        RECT 32.805 205.795 33.095 205.840 ;
        RECT 34.170 205.795 34.490 205.855 ;
        RECT 32.805 205.655 34.490 205.795 ;
        RECT 34.720 205.795 34.860 205.995 ;
        RECT 35.065 205.795 35.355 205.840 ;
        RECT 34.720 205.655 35.355 205.795 ;
        RECT 32.805 205.610 33.095 205.655 ;
        RECT 34.170 205.595 34.490 205.655 ;
        RECT 35.065 205.610 35.355 205.655 ;
        RECT 35.550 205.595 35.870 205.855 ;
        RECT 36.100 205.790 36.240 206.335 ;
        RECT 36.930 206.275 37.250 206.335 ;
        RECT 44.380 206.335 48.660 206.475 ;
        RECT 37.850 206.135 38.170 206.195 ;
        RECT 37.850 205.995 42.680 206.135 ;
        RECT 37.850 205.935 38.170 205.995 ;
        RECT 36.605 205.795 36.895 205.840 ;
        RECT 38.310 205.795 38.630 205.855 ;
        RECT 25.905 205.315 29.340 205.455 ;
        RECT 30.045 205.455 30.335 205.500 ;
        RECT 35.640 205.455 35.780 205.595 ;
        RECT 36.025 205.560 36.315 205.790 ;
        RECT 36.605 205.655 38.630 205.795 ;
        RECT 36.605 205.610 36.895 205.655 ;
        RECT 38.310 205.595 38.630 205.655 ;
        RECT 38.785 205.795 39.075 205.840 ;
        RECT 39.690 205.795 40.010 205.855 ;
        RECT 38.785 205.655 40.010 205.795 ;
        RECT 38.785 205.610 39.075 205.655 ;
        RECT 39.690 205.595 40.010 205.655 ;
        RECT 40.150 205.795 40.470 205.855 ;
        RECT 42.540 205.840 42.680 205.995 ;
        RECT 44.380 205.840 44.520 206.335 ;
        RECT 40.625 205.795 40.915 205.840 ;
        RECT 40.150 205.655 40.915 205.795 ;
        RECT 40.150 205.595 40.470 205.655 ;
        RECT 40.625 205.610 40.915 205.655 ;
        RECT 42.465 205.610 42.755 205.840 ;
        RECT 44.305 205.610 44.595 205.840 ;
        RECT 46.590 205.595 46.910 205.855 ;
        RECT 47.525 205.610 47.815 205.840 ;
        RECT 30.045 205.315 35.780 205.455 ;
        RECT 25.905 205.270 26.195 205.315 ;
        RECT 30.045 205.270 30.335 205.315 ;
        RECT 37.850 205.255 38.170 205.515 ;
        RECT 39.780 205.455 39.920 205.595 ;
        RECT 41.085 205.455 41.375 205.500 ;
        RECT 42.925 205.455 43.215 205.500 ;
        RECT 39.780 205.315 40.840 205.455 ;
        RECT 21.750 205.115 22.070 205.175 ;
        RECT 16.780 204.975 22.070 205.115 ;
        RECT 21.750 204.915 22.070 204.975 ;
        RECT 22.670 205.115 22.990 205.175 ;
        RECT 40.165 205.115 40.455 205.160 ;
        RECT 22.670 204.975 40.455 205.115 ;
        RECT 40.700 205.115 40.840 205.315 ;
        RECT 41.085 205.315 43.215 205.455 ;
        RECT 41.085 205.270 41.375 205.315 ;
        RECT 42.925 205.270 43.215 205.315 ;
        RECT 43.830 205.255 44.150 205.515 ;
        RECT 44.765 205.270 45.055 205.500 ;
        RECT 45.225 205.455 45.515 205.500 ;
        RECT 47.050 205.455 47.370 205.515 ;
        RECT 45.225 205.315 47.370 205.455 ;
        RECT 47.600 205.455 47.740 205.610 ;
        RECT 47.970 205.595 48.290 205.855 ;
        RECT 48.520 205.840 48.660 206.335 ;
        RECT 49.810 206.275 50.130 206.535 ;
        RECT 52.125 206.290 52.415 206.520 ;
        RECT 48.890 206.135 49.210 206.195 ;
        RECT 49.900 206.135 50.040 206.275 ;
        RECT 52.200 206.135 52.340 206.290 ;
        RECT 57.630 206.275 57.950 206.535 ;
        RECT 58.090 206.275 58.410 206.535 ;
        RECT 60.850 206.475 61.170 206.535 ;
        RECT 76.490 206.475 76.810 206.535 ;
        RECT 60.850 206.335 76.810 206.475 ;
        RECT 60.850 206.275 61.170 206.335 ;
        RECT 76.490 206.275 76.810 206.335 ;
        RECT 78.790 206.475 79.110 206.535 ;
        RECT 83.850 206.475 84.170 206.535 ;
        RECT 99.030 206.475 99.350 206.535 ;
        RECT 100.425 206.475 100.715 206.520 ;
        RECT 78.790 206.335 99.350 206.475 ;
        RECT 78.790 206.275 79.110 206.335 ;
        RECT 83.850 206.275 84.170 206.335 ;
        RECT 99.030 206.275 99.350 206.335 ;
        RECT 99.580 206.335 100.715 206.475 ;
        RECT 55.805 206.135 56.095 206.180 ;
        RECT 58.550 206.135 58.870 206.195 ;
        RECT 61.770 206.135 62.090 206.195 ;
        RECT 48.890 205.995 51.420 206.135 ;
        RECT 52.200 205.995 55.105 206.135 ;
        RECT 48.890 205.935 49.210 205.995 ;
        RECT 48.445 205.795 48.735 205.840 ;
        RECT 49.350 205.795 49.670 205.855 ;
        RECT 48.445 205.655 49.670 205.795 ;
        RECT 48.445 205.610 48.735 205.655 ;
        RECT 49.350 205.595 49.670 205.655 ;
        RECT 49.810 205.795 50.130 205.855 ;
        RECT 51.280 205.840 51.420 205.995 ;
        RECT 50.285 205.795 50.575 205.840 ;
        RECT 49.810 205.655 50.575 205.795 ;
        RECT 49.810 205.595 50.130 205.655 ;
        RECT 50.285 205.610 50.575 205.655 ;
        RECT 51.205 205.610 51.495 205.840 ;
        RECT 53.490 205.795 53.810 205.855 ;
        RECT 53.290 205.655 53.810 205.795 ;
        RECT 53.490 205.595 53.810 205.655 ;
        RECT 53.950 205.595 54.270 205.855 ;
        RECT 54.410 205.595 54.730 205.855 ;
        RECT 54.965 205.840 55.105 205.995 ;
        RECT 55.805 205.995 58.870 206.135 ;
        RECT 55.805 205.950 56.095 205.995 ;
        RECT 58.550 205.935 58.870 205.995 ;
        RECT 59.100 205.995 62.090 206.135 ;
        RECT 54.890 205.610 55.180 205.840 ;
        RECT 56.250 205.595 56.570 205.855 ;
        RECT 59.100 205.840 59.240 205.995 ;
        RECT 61.770 205.935 62.090 205.995 ;
        RECT 64.545 206.135 64.835 206.180 ;
        RECT 65.450 206.135 65.770 206.195 ;
        RECT 64.545 205.995 65.770 206.135 ;
        RECT 64.545 205.950 64.835 205.995 ;
        RECT 65.450 205.935 65.770 205.995 ;
        RECT 67.750 205.935 68.070 206.195 ;
        RECT 69.590 206.135 69.910 206.195 ;
        RECT 70.525 206.135 70.815 206.180 ;
        RECT 71.445 206.135 71.735 206.180 ;
        RECT 74.190 206.135 74.510 206.195 ;
        RECT 69.590 205.995 70.815 206.135 ;
        RECT 69.590 205.935 69.910 205.995 ;
        RECT 70.525 205.950 70.815 205.995 ;
        RECT 71.060 205.995 71.735 206.135 ;
        RECT 56.750 205.610 57.040 205.840 ;
        RECT 59.025 205.610 59.315 205.840 ;
        RECT 59.485 205.610 59.775 205.840 ;
        RECT 59.945 205.610 60.235 205.840 ;
        RECT 60.865 205.795 61.155 205.840 ;
        RECT 62.230 205.795 62.550 205.855 ;
        RECT 60.865 205.655 62.550 205.795 ;
        RECT 60.865 205.610 61.155 205.655 ;
        RECT 53.575 205.455 53.715 205.595 ;
        RECT 56.825 205.455 56.965 205.610 ;
        RECT 47.600 205.315 56.965 205.455 ;
        RECT 57.170 205.455 57.490 205.515 ;
        RECT 59.560 205.455 59.700 205.610 ;
        RECT 57.170 205.315 59.700 205.455 ;
        RECT 60.020 205.455 60.160 205.610 ;
        RECT 62.230 205.595 62.550 205.655 ;
        RECT 62.705 205.795 62.995 205.840 ;
        RECT 63.150 205.795 63.470 205.855 ;
        RECT 62.705 205.655 63.470 205.795 ;
        RECT 62.705 205.610 62.995 205.655 ;
        RECT 63.150 205.595 63.470 205.655 ;
        RECT 64.070 205.595 64.390 205.855 ;
        RECT 64.990 205.795 65.310 205.855 ;
        RECT 64.990 205.655 69.360 205.795 ;
        RECT 64.990 205.595 65.310 205.655 ;
        RECT 61.310 205.455 61.630 205.515 ;
        RECT 60.020 205.315 61.630 205.455 ;
        RECT 45.225 205.270 45.515 205.315 ;
        RECT 44.840 205.115 44.980 205.270 ;
        RECT 47.050 205.255 47.370 205.315 ;
        RECT 57.170 205.255 57.490 205.315 ;
        RECT 61.310 205.255 61.630 205.315 ;
        RECT 61.785 205.270 62.075 205.500 ;
        RECT 63.625 205.455 63.915 205.500 ;
        RECT 68.225 205.455 68.515 205.500 ;
        RECT 63.625 205.315 68.515 205.455 ;
        RECT 63.625 205.270 63.915 205.315 ;
        RECT 68.225 205.270 68.515 205.315 ;
        RECT 47.970 205.115 48.290 205.175 ;
        RECT 40.700 204.975 48.290 205.115 ;
        RECT 22.670 204.915 22.990 204.975 ;
        RECT 40.165 204.930 40.455 204.975 ;
        RECT 47.970 204.915 48.290 204.975 ;
        RECT 51.650 205.115 51.970 205.175 ;
        RECT 58.090 205.115 58.410 205.175 ;
        RECT 51.650 204.975 58.410 205.115 ;
        RECT 51.650 204.915 51.970 204.975 ;
        RECT 58.090 204.915 58.410 204.975 ;
        RECT 59.470 205.115 59.790 205.175 ;
        RECT 61.860 205.115 62.000 205.270 ;
        RECT 68.670 205.255 68.990 205.515 ;
        RECT 64.990 205.115 65.310 205.175 ;
        RECT 59.470 204.975 65.310 205.115 ;
        RECT 59.470 204.915 59.790 204.975 ;
        RECT 64.990 204.915 65.310 204.975 ;
        RECT 65.925 205.115 66.215 205.160 ;
        RECT 66.370 205.115 66.690 205.175 ;
        RECT 65.925 204.975 66.690 205.115 ;
        RECT 69.220 205.115 69.360 205.655 ;
        RECT 70.050 205.595 70.370 205.855 ;
        RECT 71.060 205.840 71.200 205.995 ;
        RECT 71.445 205.950 71.735 205.995 ;
        RECT 73.360 205.995 74.510 206.135 ;
        RECT 70.985 205.610 71.275 205.840 ;
        RECT 71.905 205.795 72.195 205.840 ;
        RECT 73.360 205.795 73.500 205.995 ;
        RECT 74.190 205.935 74.510 205.995 ;
        RECT 79.250 206.135 79.570 206.195 ;
        RECT 82.945 206.135 83.235 206.180 ;
        RECT 84.310 206.135 84.630 206.195 ;
        RECT 79.250 205.995 82.240 206.135 ;
        RECT 79.250 205.935 79.570 205.995 ;
        RECT 82.100 205.855 82.240 205.995 ;
        RECT 82.945 205.995 84.630 206.135 ;
        RECT 82.945 205.950 83.235 205.995 ;
        RECT 84.310 205.935 84.630 205.995 ;
        RECT 87.530 206.135 87.850 206.195 ;
        RECT 91.210 206.135 91.530 206.195 ;
        RECT 92.145 206.135 92.435 206.180 ;
        RECT 99.580 206.135 99.720 206.335 ;
        RECT 100.425 206.290 100.715 206.335 ;
        RECT 102.710 206.475 103.030 206.535 ;
        RECT 108.230 206.475 108.550 206.535 ;
        RECT 102.710 206.335 108.550 206.475 ;
        RECT 102.710 206.275 103.030 206.335 ;
        RECT 108.230 206.275 108.550 206.335 ;
        RECT 109.150 206.475 109.470 206.535 ;
        RECT 109.625 206.475 109.915 206.520 ;
        RECT 109.150 206.335 109.915 206.475 ;
        RECT 109.150 206.275 109.470 206.335 ;
        RECT 109.625 206.290 109.915 206.335 ;
        RECT 111.925 206.475 112.215 206.520 ;
        RECT 119.730 206.475 120.050 206.535 ;
        RECT 111.925 206.335 120.050 206.475 ;
        RECT 111.925 206.290 112.215 206.335 ;
        RECT 119.730 206.275 120.050 206.335 ;
        RECT 120.650 206.475 120.970 206.535 ;
        RECT 121.125 206.475 121.415 206.520 ;
        RECT 120.650 206.335 121.415 206.475 ;
        RECT 120.650 206.275 120.970 206.335 ;
        RECT 121.125 206.290 121.415 206.335 ;
        RECT 129.390 206.275 129.710 206.535 ;
        RECT 129.850 206.475 130.170 206.535 ;
        RECT 137.210 206.475 137.530 206.535 ;
        RECT 129.850 206.335 137.530 206.475 ;
        RECT 129.850 206.275 130.170 206.335 ;
        RECT 137.210 206.275 137.530 206.335 ;
        RECT 145.490 206.275 145.810 206.535 ;
        RECT 105.470 206.135 105.790 206.195 ;
        RECT 87.530 205.995 92.435 206.135 ;
        RECT 87.530 205.935 87.850 205.995 ;
        RECT 91.210 205.935 91.530 205.995 ;
        RECT 92.145 205.950 92.435 205.995 ;
        RECT 94.980 205.995 99.720 206.135 ;
        RECT 102.800 205.995 105.790 206.135 ;
        RECT 71.905 205.655 73.500 205.795 ;
        RECT 73.745 205.795 74.035 205.840 ;
        RECT 81.550 205.795 81.870 205.855 ;
        RECT 73.745 205.655 81.870 205.795 ;
        RECT 71.905 205.610 72.195 205.655 ;
        RECT 73.745 205.610 74.035 205.655 ;
        RECT 71.430 205.455 71.750 205.515 ;
        RECT 71.980 205.455 72.120 205.610 ;
        RECT 81.550 205.595 81.870 205.655 ;
        RECT 82.010 205.795 82.330 205.855 ;
        RECT 85.705 205.795 85.995 205.840 ;
        RECT 82.010 205.655 85.995 205.795 ;
        RECT 82.010 205.595 82.330 205.655 ;
        RECT 85.705 205.610 85.995 205.655 ;
        RECT 86.150 205.595 86.470 205.855 ;
        RECT 86.610 205.595 86.930 205.855 ;
        RECT 87.085 205.795 87.375 205.840 ;
        RECT 92.590 205.795 92.910 205.855 ;
        RECT 94.430 205.795 94.750 205.855 ;
        RECT 94.980 205.840 95.120 205.995 ;
        RECT 87.085 205.655 92.360 205.795 ;
        RECT 87.085 205.610 87.375 205.655 ;
        RECT 71.430 205.315 72.120 205.455 ;
        RECT 72.350 205.455 72.670 205.515 ;
        RECT 78.790 205.455 79.110 205.515 ;
        RECT 72.350 205.315 79.110 205.455 ;
        RECT 71.430 205.255 71.750 205.315 ;
        RECT 72.350 205.255 72.670 205.315 ;
        RECT 78.790 205.255 79.110 205.315 ;
        RECT 80.630 205.455 80.950 205.515 ;
        RECT 83.405 205.455 83.695 205.500 ;
        RECT 86.700 205.455 86.840 205.595 ;
        RECT 80.630 205.315 83.695 205.455 ;
        RECT 80.630 205.255 80.950 205.315 ;
        RECT 83.405 205.270 83.695 205.315 ;
        RECT 85.780 205.315 86.840 205.455 ;
        RECT 87.990 205.455 88.310 205.515 ;
        RECT 88.465 205.455 88.755 205.500 ;
        RECT 87.990 205.315 88.755 205.455 ;
        RECT 85.780 205.175 85.920 205.315 ;
        RECT 87.990 205.255 88.310 205.315 ;
        RECT 88.465 205.270 88.755 205.315 ;
        RECT 90.750 205.255 91.070 205.515 ;
        RECT 92.220 205.455 92.360 205.655 ;
        RECT 92.590 205.655 94.750 205.795 ;
        RECT 92.590 205.595 92.910 205.655 ;
        RECT 94.430 205.595 94.750 205.655 ;
        RECT 94.905 205.610 95.195 205.840 ;
        RECT 95.825 205.795 96.115 205.840 ;
        RECT 96.730 205.795 97.050 205.855 ;
        RECT 98.125 205.795 98.415 205.840 ;
        RECT 95.825 205.655 96.500 205.795 ;
        RECT 95.825 205.610 96.115 205.655 ;
        RECT 92.220 205.315 96.040 205.455 ;
        RECT 84.325 205.115 84.615 205.160 ;
        RECT 85.690 205.115 86.010 205.175 ;
        RECT 69.220 204.975 73.500 205.115 ;
        RECT 65.925 204.930 66.215 204.975 ;
        RECT 66.370 204.915 66.690 204.975 ;
        RECT 14.060 204.775 14.380 204.835 ;
        RECT 17.625 204.775 17.915 204.820 ;
        RECT 14.060 204.635 17.915 204.775 ;
        RECT 14.060 204.575 14.380 204.635 ;
        RECT 17.625 204.590 17.915 204.635 ;
        RECT 18.530 204.775 18.850 204.835 ;
        RECT 19.005 204.775 19.295 204.820 ;
        RECT 18.530 204.635 19.295 204.775 ;
        RECT 18.530 204.575 18.850 204.635 ;
        RECT 19.005 204.590 19.295 204.635 ;
        RECT 24.970 204.775 25.290 204.835 ;
        RECT 25.445 204.775 25.735 204.820 ;
        RECT 24.970 204.635 25.735 204.775 ;
        RECT 24.970 204.575 25.290 204.635 ;
        RECT 25.445 204.590 25.735 204.635 ;
        RECT 27.730 204.575 28.050 204.835 ;
        RECT 30.490 204.575 30.810 204.835 ;
        RECT 30.950 204.775 31.270 204.835 ;
        RECT 31.425 204.775 31.715 204.820 ;
        RECT 30.950 204.635 31.715 204.775 ;
        RECT 30.950 204.575 31.270 204.635 ;
        RECT 31.425 204.590 31.715 204.635 ;
        RECT 31.870 204.775 32.190 204.835 ;
        RECT 32.345 204.775 32.635 204.820 ;
        RECT 31.870 204.635 32.635 204.775 ;
        RECT 31.870 204.575 32.190 204.635 ;
        RECT 32.345 204.590 32.635 204.635 ;
        RECT 34.630 204.775 34.950 204.835 ;
        RECT 35.565 204.775 35.855 204.820 ;
        RECT 34.630 204.635 35.855 204.775 ;
        RECT 34.630 204.575 34.950 204.635 ;
        RECT 35.565 204.590 35.855 204.635 ;
        RECT 36.930 204.575 37.250 204.835 ;
        RECT 42.005 204.775 42.295 204.820 ;
        RECT 49.350 204.775 49.670 204.835 ;
        RECT 42.005 204.635 49.670 204.775 ;
        RECT 42.005 204.590 42.295 204.635 ;
        RECT 49.350 204.575 49.670 204.635 ;
        RECT 50.730 204.775 51.050 204.835 ;
        RECT 53.950 204.775 54.270 204.835 ;
        RECT 50.730 204.635 54.270 204.775 ;
        RECT 50.730 204.575 51.050 204.635 ;
        RECT 53.950 204.575 54.270 204.635 ;
        RECT 67.290 204.775 67.610 204.835 ;
        RECT 71.890 204.775 72.210 204.835 ;
        RECT 73.360 204.820 73.500 204.975 ;
        RECT 84.325 204.975 86.010 205.115 ;
        RECT 84.325 204.930 84.615 204.975 ;
        RECT 85.690 204.915 86.010 204.975 ;
        RECT 86.610 204.915 86.930 205.175 ;
        RECT 89.385 204.930 89.675 205.160 ;
        RECT 90.290 205.115 90.610 205.175 ;
        RECT 95.365 205.115 95.655 205.160 ;
        RECT 90.290 204.975 95.655 205.115 ;
        RECT 67.290 204.635 72.210 204.775 ;
        RECT 67.290 204.575 67.610 204.635 ;
        RECT 71.890 204.575 72.210 204.635 ;
        RECT 73.285 204.775 73.575 204.820 ;
        RECT 76.030 204.775 76.350 204.835 ;
        RECT 73.285 204.635 76.350 204.775 ;
        RECT 73.285 204.590 73.575 204.635 ;
        RECT 76.030 204.575 76.350 204.635 ;
        RECT 83.850 204.775 84.170 204.835 ;
        RECT 88.910 204.775 89.230 204.835 ;
        RECT 83.850 204.635 89.230 204.775 ;
        RECT 89.460 204.775 89.600 204.930 ;
        RECT 90.290 204.915 90.610 204.975 ;
        RECT 95.365 204.930 95.655 204.975 ;
        RECT 92.590 204.775 92.910 204.835 ;
        RECT 89.460 204.635 92.910 204.775 ;
        RECT 95.900 204.775 96.040 205.315 ;
        RECT 96.360 205.160 96.500 205.655 ;
        RECT 96.730 205.655 98.415 205.795 ;
        RECT 100.870 205.785 101.190 205.855 ;
        RECT 102.800 205.840 102.940 205.995 ;
        RECT 105.470 205.935 105.790 205.995 ;
        RECT 105.930 205.935 106.250 206.195 ;
        RECT 120.190 206.135 120.510 206.195 ;
        RECT 110.620 205.995 120.510 206.135 ;
        RECT 96.730 205.595 97.050 205.655 ;
        RECT 98.125 205.610 98.415 205.655 ;
        RECT 100.500 205.645 101.190 205.785 ;
        RECT 98.570 205.255 98.890 205.515 ;
        RECT 99.045 205.270 99.335 205.500 ;
        RECT 100.500 205.455 100.640 205.645 ;
        RECT 100.870 205.595 101.190 205.645 ;
        RECT 102.725 205.610 103.015 205.840 ;
        RECT 104.090 205.595 104.410 205.855 ;
        RECT 104.550 205.595 104.870 205.855 ;
        RECT 110.620 205.840 110.760 205.995 ;
        RECT 120.190 205.935 120.510 205.995 ;
        RECT 121.570 206.135 121.890 206.195 ;
        RECT 125.725 206.135 126.015 206.180 ;
        RECT 126.170 206.135 126.490 206.195 ;
        RECT 128.470 206.135 128.790 206.195 ;
        RECT 134.465 206.135 134.755 206.180 ;
        RECT 121.570 205.995 126.490 206.135 ;
        RECT 121.570 205.935 121.890 205.995 ;
        RECT 125.725 205.950 126.015 205.995 ;
        RECT 126.170 205.935 126.490 205.995 ;
        RECT 127.180 205.995 128.790 206.135 ;
        RECT 105.025 205.610 105.315 205.840 ;
        RECT 110.545 205.610 110.835 205.840 ;
        RECT 101.345 205.455 101.635 205.500 ;
        RECT 100.500 205.315 101.635 205.455 ;
        RECT 101.345 205.270 101.635 205.315 ;
        RECT 101.805 205.270 102.095 205.500 ;
        RECT 102.265 205.455 102.555 205.500 ;
        RECT 102.265 205.315 102.940 205.455 ;
        RECT 102.265 205.270 102.555 205.315 ;
        RECT 96.285 204.930 96.575 205.160 ;
        RECT 97.650 205.115 97.970 205.175 ;
        RECT 99.120 205.115 99.260 205.270 ;
        RECT 97.650 204.975 99.260 205.115 ;
        RECT 99.490 205.115 99.810 205.175 ;
        RECT 101.880 205.115 102.020 205.270 ;
        RECT 99.490 204.975 102.020 205.115 ;
        RECT 102.800 205.115 102.940 205.315 ;
        RECT 104.640 205.115 104.780 205.595 ;
        RECT 105.100 205.175 105.240 205.610 ;
        RECT 112.830 205.595 113.150 205.855 ;
        RECT 114.210 205.595 114.530 205.855 ;
        RECT 116.510 205.795 116.830 205.855 ;
        RECT 117.445 205.795 117.735 205.840 ;
        RECT 119.745 205.795 120.035 205.840 ;
        RECT 122.030 205.795 122.350 205.855 ;
        RECT 116.065 205.560 116.355 205.790 ;
        RECT 116.510 205.655 117.735 205.795 ;
        RECT 116.510 205.595 116.830 205.655 ;
        RECT 117.445 205.610 117.735 205.655 ;
        RECT 117.980 205.655 122.350 205.795 ;
        RECT 106.865 205.455 107.155 205.500 ;
        RECT 107.310 205.455 107.630 205.515 ;
        RECT 106.865 205.315 107.630 205.455 ;
        RECT 106.865 205.270 107.155 205.315 ;
        RECT 107.310 205.255 107.630 205.315 ;
        RECT 110.990 205.255 111.310 205.515 ;
        RECT 112.385 205.455 112.675 205.500 ;
        RECT 115.590 205.455 115.910 205.515 ;
        RECT 112.385 205.315 115.910 205.455 ;
        RECT 112.385 205.270 112.675 205.315 ;
        RECT 115.590 205.255 115.910 205.315 ;
        RECT 102.800 204.975 104.780 205.115 ;
        RECT 105.010 205.115 105.330 205.175 ;
        RECT 107.770 205.115 108.090 205.175 ;
        RECT 108.245 205.115 108.535 205.160 ;
        RECT 105.010 204.975 108.535 205.115 ;
        RECT 97.650 204.915 97.970 204.975 ;
        RECT 99.490 204.915 99.810 204.975 ;
        RECT 105.010 204.915 105.330 204.975 ;
        RECT 107.770 204.915 108.090 204.975 ;
        RECT 108.245 204.930 108.535 204.975 ;
        RECT 109.165 205.115 109.455 205.160 ;
        RECT 116.140 205.115 116.280 205.560 ;
        RECT 116.970 205.455 117.290 205.515 ;
        RECT 117.980 205.455 118.120 205.655 ;
        RECT 119.745 205.610 120.035 205.655 ;
        RECT 122.030 205.595 122.350 205.655 ;
        RECT 123.410 205.795 123.730 205.855 ;
        RECT 123.885 205.795 124.175 205.840 ;
        RECT 123.410 205.655 124.175 205.795 ;
        RECT 123.410 205.595 123.730 205.655 ;
        RECT 123.885 205.610 124.175 205.655 ;
        RECT 124.805 205.795 125.095 205.840 ;
        RECT 125.250 205.795 125.570 205.855 ;
        RECT 127.180 205.840 127.320 205.995 ;
        RECT 128.470 205.935 128.790 205.995 ;
        RECT 129.020 205.995 134.755 206.135 ;
        RECT 129.020 205.855 129.160 205.995 ;
        RECT 134.465 205.950 134.755 205.995 ;
        RECT 124.805 205.655 125.570 205.795 ;
        RECT 124.805 205.610 125.095 205.655 ;
        RECT 125.250 205.595 125.570 205.655 ;
        RECT 127.105 205.610 127.395 205.840 ;
        RECT 127.550 205.595 127.870 205.855 ;
        RECT 128.930 205.595 129.250 205.855 ;
        RECT 129.850 205.595 130.170 205.855 ;
        RECT 130.310 205.595 130.630 205.855 ;
        RECT 131.230 205.595 131.550 205.855 ;
        RECT 132.625 205.610 132.915 205.840 ;
        RECT 137.685 205.795 137.975 205.840 ;
        RECT 139.050 205.795 139.370 205.855 ;
        RECT 137.685 205.655 139.370 205.795 ;
        RECT 137.685 205.610 137.975 205.655 ;
        RECT 116.970 205.315 118.120 205.455 ;
        RECT 118.825 205.455 119.115 205.500 ;
        RECT 128.470 205.455 128.790 205.515 ;
        RECT 132.700 205.455 132.840 205.610 ;
        RECT 139.050 205.595 139.370 205.655 ;
        RECT 140.890 205.595 141.210 205.855 ;
        RECT 144.110 205.795 144.430 205.855 ;
        RECT 144.585 205.795 144.875 205.840 ;
        RECT 144.110 205.655 144.875 205.795 ;
        RECT 144.110 205.595 144.430 205.655 ;
        RECT 144.585 205.610 144.875 205.655 ;
        RECT 133.530 205.455 133.850 205.515 ;
        RECT 118.825 205.315 122.720 205.455 ;
        RECT 116.970 205.255 117.290 205.315 ;
        RECT 118.825 205.270 119.115 205.315 ;
        RECT 117.430 205.115 117.750 205.175 ;
        RECT 109.165 204.975 117.750 205.115 ;
        RECT 109.165 204.930 109.455 204.975 ;
        RECT 117.430 204.915 117.750 204.975 ;
        RECT 103.630 204.775 103.950 204.835 ;
        RECT 95.900 204.635 103.950 204.775 ;
        RECT 83.850 204.575 84.170 204.635 ;
        RECT 88.910 204.575 89.230 204.635 ;
        RECT 92.590 204.575 92.910 204.635 ;
        RECT 103.630 204.575 103.950 204.635 ;
        RECT 113.290 204.575 113.610 204.835 ;
        RECT 115.605 204.775 115.895 204.820 ;
        RECT 118.900 204.775 119.040 205.270 ;
        RECT 119.270 205.115 119.590 205.175 ;
        RECT 122.580 205.115 122.720 205.315 ;
        RECT 128.470 205.315 133.850 205.455 ;
        RECT 128.470 205.255 128.790 205.315 ;
        RECT 133.530 205.255 133.850 205.315 ;
        RECT 132.150 205.115 132.470 205.175 ;
        RECT 119.270 204.975 122.260 205.115 ;
        RECT 122.580 204.975 132.470 205.115 ;
        RECT 119.270 204.915 119.590 204.975 ;
        RECT 115.605 204.635 119.040 204.775 ;
        RECT 115.605 204.590 115.895 204.635 ;
        RECT 119.730 204.575 120.050 204.835 ;
        RECT 120.665 204.775 120.955 204.820 ;
        RECT 121.110 204.775 121.430 204.835 ;
        RECT 122.120 204.820 122.260 204.975 ;
        RECT 132.150 204.915 132.470 204.975 ;
        RECT 132.610 205.115 132.930 205.175 ;
        RECT 132.610 204.975 133.760 205.115 ;
        RECT 132.610 204.915 132.930 204.975 ;
        RECT 120.665 204.635 121.430 204.775 ;
        RECT 120.665 204.590 120.955 204.635 ;
        RECT 121.110 204.575 121.430 204.635 ;
        RECT 122.045 204.590 122.335 204.820 ;
        RECT 124.330 204.775 124.650 204.835 ;
        RECT 128.025 204.775 128.315 204.820 ;
        RECT 124.330 204.635 128.315 204.775 ;
        RECT 124.330 204.575 124.650 204.635 ;
        RECT 128.025 204.590 128.315 204.635 ;
        RECT 131.245 204.775 131.535 204.820 ;
        RECT 133.070 204.775 133.390 204.835 ;
        RECT 133.620 204.820 133.760 204.975 ;
        RECT 131.245 204.635 133.390 204.775 ;
        RECT 131.245 204.590 131.535 204.635 ;
        RECT 133.070 204.575 133.390 204.635 ;
        RECT 133.545 204.590 133.835 204.820 ;
        RECT 141.810 204.575 142.130 204.835 ;
        RECT 13.860 203.955 147.720 204.435 ;
        RECT 18.940 203.755 19.230 203.800 ;
        RECT 27.285 203.755 27.575 203.800 ;
        RECT 18.940 203.615 27.575 203.755 ;
        RECT 18.940 203.570 19.230 203.615 ;
        RECT 27.285 203.570 27.575 203.615 ;
        RECT 32.805 203.755 33.095 203.800 ;
        RECT 34.170 203.755 34.490 203.815 ;
        RECT 32.805 203.615 34.490 203.755 ;
        RECT 32.805 203.570 33.095 203.615 ;
        RECT 34.170 203.555 34.490 203.615 ;
        RECT 36.470 203.555 36.790 203.815 ;
        RECT 36.930 203.755 37.250 203.815 ;
        RECT 45.210 203.755 45.530 203.815 ;
        RECT 66.370 203.755 66.690 203.815 ;
        RECT 36.930 203.615 66.690 203.755 ;
        RECT 36.930 203.555 37.250 203.615 ;
        RECT 45.210 203.555 45.530 203.615 ;
        RECT 66.370 203.555 66.690 203.615 ;
        RECT 66.830 203.755 67.150 203.815 ;
        RECT 67.305 203.755 67.595 203.800 ;
        RECT 66.830 203.615 67.595 203.755 ;
        RECT 66.830 203.555 67.150 203.615 ;
        RECT 67.305 203.570 67.595 203.615 ;
        RECT 70.970 203.555 71.290 203.815 ;
        RECT 73.285 203.570 73.575 203.800 ;
        RECT 75.125 203.755 75.415 203.800 ;
        RECT 76.950 203.755 77.270 203.815 ;
        RECT 75.125 203.615 77.270 203.755 ;
        RECT 75.125 203.570 75.415 203.615 ;
        RECT 13.930 203.415 14.250 203.475 ;
        RECT 15.785 203.415 16.075 203.460 ;
        RECT 13.930 203.275 16.075 203.415 ;
        RECT 13.930 203.215 14.250 203.275 ;
        RECT 15.785 203.230 16.075 203.275 ;
        RECT 18.495 203.415 18.785 203.460 ;
        RECT 20.385 203.415 20.675 203.460 ;
        RECT 23.505 203.415 23.795 203.460 ;
        RECT 18.495 203.275 23.795 203.415 ;
        RECT 18.495 203.230 18.785 203.275 ;
        RECT 20.385 203.230 20.675 203.275 ;
        RECT 23.505 203.230 23.795 203.275 ;
        RECT 26.365 203.415 26.655 203.460 ;
        RECT 31.410 203.415 31.730 203.475 ;
        RECT 33.265 203.415 33.555 203.460 ;
        RECT 26.365 203.275 33.555 203.415 ;
        RECT 26.365 203.230 26.655 203.275 ;
        RECT 31.410 203.215 31.730 203.275 ;
        RECT 33.265 203.230 33.555 203.275 ;
        RECT 37.390 203.415 37.710 203.475 ;
        RECT 50.285 203.415 50.575 203.460 ;
        RECT 37.390 203.275 50.575 203.415 ;
        RECT 37.390 203.215 37.710 203.275 ;
        RECT 50.285 203.230 50.575 203.275 ;
        RECT 50.730 203.415 51.050 203.475 ;
        RECT 54.410 203.415 54.730 203.475 ;
        RECT 50.730 203.275 54.730 203.415 ;
        RECT 50.730 203.215 51.050 203.275 ;
        RECT 54.410 203.215 54.730 203.275 ;
        RECT 54.885 203.415 55.175 203.460 ;
        RECT 55.790 203.415 56.110 203.475 ;
        RECT 54.885 203.275 56.110 203.415 ;
        RECT 54.885 203.230 55.175 203.275 ;
        RECT 55.790 203.215 56.110 203.275 ;
        RECT 56.725 203.415 57.015 203.460 ;
        RECT 64.070 203.415 64.390 203.475 ;
        RECT 56.725 203.275 64.390 203.415 ;
        RECT 56.725 203.230 57.015 203.275 ;
        RECT 64.070 203.215 64.390 203.275 ;
        RECT 65.910 203.415 66.230 203.475 ;
        RECT 73.360 203.415 73.500 203.570 ;
        RECT 76.950 203.555 77.270 203.615 ;
        RECT 81.550 203.755 81.870 203.815 ;
        RECT 85.245 203.755 85.535 203.800 ;
        RECT 87.990 203.755 88.310 203.815 ;
        RECT 106.850 203.755 107.170 203.815 ;
        RECT 81.550 203.615 85.535 203.755 ;
        RECT 81.550 203.555 81.870 203.615 ;
        RECT 85.245 203.570 85.535 203.615 ;
        RECT 85.780 203.615 88.310 203.755 ;
        RECT 85.780 203.415 85.920 203.615 ;
        RECT 87.990 203.555 88.310 203.615 ;
        RECT 88.540 203.615 107.170 203.755 ;
        RECT 65.910 203.275 73.500 203.415 ;
        RECT 77.040 203.275 85.920 203.415 ;
        RECT 65.910 203.215 66.230 203.275 ;
        RECT 17.625 203.075 17.915 203.120 ;
        RECT 18.990 203.075 19.310 203.135 ;
        RECT 17.625 202.935 19.310 203.075 ;
        RECT 17.625 202.890 17.915 202.935 ;
        RECT 18.990 202.875 19.310 202.935 ;
        RECT 21.750 203.075 22.070 203.135 ;
        RECT 30.505 203.075 30.795 203.120 ;
        RECT 35.090 203.075 35.410 203.135 ;
        RECT 66.370 203.075 66.690 203.135 ;
        RECT 21.750 202.935 29.800 203.075 ;
        RECT 21.750 202.875 22.070 202.935 ;
        RECT 16.690 202.535 17.010 202.795 ;
        RECT 18.090 202.735 18.380 202.780 ;
        RECT 19.925 202.735 20.215 202.780 ;
        RECT 23.505 202.735 23.795 202.780 ;
        RECT 18.090 202.595 23.795 202.735 ;
        RECT 18.090 202.550 18.380 202.595 ;
        RECT 19.925 202.550 20.215 202.595 ;
        RECT 23.505 202.550 23.795 202.595 ;
        RECT 24.585 202.440 24.875 202.755 ;
        RECT 27.730 202.735 28.050 202.795 ;
        RECT 29.125 202.735 29.415 202.780 ;
        RECT 27.730 202.595 29.415 202.735 ;
        RECT 27.730 202.535 28.050 202.595 ;
        RECT 29.125 202.550 29.415 202.595 ;
        RECT 21.285 202.395 21.935 202.440 ;
        RECT 24.585 202.395 25.175 202.440 ;
        RECT 26.350 202.395 26.670 202.455 ;
        RECT 21.285 202.255 26.670 202.395 ;
        RECT 29.660 202.395 29.800 202.935 ;
        RECT 30.505 202.935 35.410 203.075 ;
        RECT 30.505 202.890 30.795 202.935 ;
        RECT 35.090 202.875 35.410 202.935 ;
        RECT 43.000 202.935 61.080 203.075 ;
        RECT 30.030 202.735 30.350 202.795 ;
        RECT 31.885 202.735 32.175 202.780 ;
        RECT 30.030 202.595 32.175 202.735 ;
        RECT 30.030 202.535 30.350 202.595 ;
        RECT 31.885 202.550 32.175 202.595 ;
        RECT 32.345 202.735 32.635 202.780 ;
        RECT 32.790 202.735 33.110 202.795 ;
        RECT 32.345 202.595 33.110 202.735 ;
        RECT 32.345 202.550 32.635 202.595 ;
        RECT 32.790 202.535 33.110 202.595 ;
        RECT 33.725 202.735 34.015 202.780 ;
        RECT 39.230 202.735 39.550 202.795 ;
        RECT 43.000 202.780 43.140 202.935 ;
        RECT 60.940 202.795 61.080 202.935 ;
        RECT 66.370 202.935 69.820 203.075 ;
        RECT 66.370 202.875 66.690 202.935 ;
        RECT 33.725 202.595 39.550 202.735 ;
        RECT 33.725 202.550 34.015 202.595 ;
        RECT 39.230 202.535 39.550 202.595 ;
        RECT 42.925 202.550 43.215 202.780 ;
        RECT 43.830 202.535 44.150 202.795 ;
        RECT 45.210 202.535 45.530 202.795 ;
        RECT 46.590 202.535 46.910 202.795 ;
        RECT 47.970 202.535 48.290 202.795 ;
        RECT 48.890 202.735 49.210 202.795 ;
        RECT 49.825 202.735 50.115 202.780 ;
        RECT 48.890 202.595 50.115 202.735 ;
        RECT 48.890 202.535 49.210 202.595 ;
        RECT 49.825 202.550 50.115 202.595 ;
        RECT 50.285 202.735 50.575 202.780 ;
        RECT 50.730 202.735 51.050 202.795 ;
        RECT 50.285 202.595 51.050 202.735 ;
        RECT 50.285 202.550 50.575 202.595 ;
        RECT 50.730 202.535 51.050 202.595 ;
        RECT 51.205 202.735 51.495 202.780 ;
        RECT 56.250 202.735 56.570 202.795 ;
        RECT 51.205 202.595 56.570 202.735 ;
        RECT 51.205 202.550 51.495 202.595 ;
        RECT 56.250 202.535 56.570 202.595 ;
        RECT 56.725 202.550 57.015 202.780 ;
        RECT 40.150 202.395 40.470 202.455 ;
        RECT 29.660 202.255 40.470 202.395 ;
        RECT 43.920 202.395 44.060 202.535 ;
        RECT 46.680 202.395 46.820 202.535 ;
        RECT 43.920 202.255 46.820 202.395 ;
        RECT 21.285 202.210 21.935 202.255 ;
        RECT 24.885 202.210 25.175 202.255 ;
        RECT 26.350 202.195 26.670 202.255 ;
        RECT 40.150 202.195 40.470 202.255 ;
        RECT 48.430 202.195 48.750 202.455 ;
        RECT 49.350 202.195 49.670 202.455 ;
        RECT 53.965 202.210 54.255 202.440 ;
        RECT 55.345 202.210 55.635 202.440 ;
        RECT 56.800 202.395 56.940 202.550 ;
        RECT 57.170 202.535 57.490 202.795 ;
        RECT 58.090 202.535 58.410 202.795 ;
        RECT 58.550 202.535 58.870 202.795 ;
        RECT 59.010 202.535 59.330 202.795 ;
        RECT 60.850 202.735 61.170 202.795 ;
        RECT 60.665 202.595 61.170 202.735 ;
        RECT 60.850 202.535 61.170 202.595 ;
        RECT 61.310 202.735 61.630 202.795 ;
        RECT 67.290 202.735 67.610 202.795 ;
        RECT 61.310 202.595 67.610 202.735 ;
        RECT 61.310 202.535 61.630 202.595 ;
        RECT 67.290 202.535 67.610 202.595 ;
        RECT 69.130 202.395 69.450 202.455 ;
        RECT 56.800 202.255 69.450 202.395 ;
        RECT 69.680 202.395 69.820 202.935 ;
        RECT 71.430 202.875 71.750 203.135 ;
        RECT 71.890 203.075 72.210 203.135 ;
        RECT 77.040 203.120 77.180 203.275 ;
        RECT 87.530 203.215 87.850 203.475 ;
        RECT 73.360 203.075 74.420 203.115 ;
        RECT 76.965 203.075 77.255 203.120 ;
        RECT 71.890 202.975 77.255 203.075 ;
        RECT 71.890 202.935 73.500 202.975 ;
        RECT 74.280 202.935 77.255 202.975 ;
        RECT 71.890 202.875 72.210 202.935 ;
        RECT 76.965 202.890 77.255 202.935 ;
        RECT 77.500 202.935 79.480 203.075 ;
        RECT 70.510 202.735 70.830 202.795 ;
        RECT 72.825 202.735 73.115 202.780 ;
        RECT 70.510 202.595 73.115 202.735 ;
        RECT 70.510 202.535 70.830 202.595 ;
        RECT 72.825 202.550 73.115 202.595 ;
        RECT 73.285 202.735 73.575 202.780 ;
        RECT 73.730 202.735 74.050 202.795 ;
        RECT 73.285 202.595 74.050 202.735 ;
        RECT 73.285 202.550 73.575 202.595 ;
        RECT 73.730 202.535 74.050 202.595 ;
        RECT 74.190 202.535 74.510 202.795 ;
        RECT 75.570 202.535 75.890 202.795 ;
        RECT 76.030 202.535 76.350 202.795 ;
        RECT 76.490 202.735 76.810 202.795 ;
        RECT 77.500 202.735 77.640 202.935 ;
        RECT 76.490 202.595 77.640 202.735 ;
        RECT 76.490 202.535 76.810 202.595 ;
        RECT 78.805 202.550 79.095 202.780 ;
        RECT 78.880 202.395 79.020 202.550 ;
        RECT 69.680 202.255 79.020 202.395 ;
        RECT 79.340 202.395 79.480 202.935 ;
        RECT 83.850 202.875 84.170 203.135 ;
        RECT 84.770 203.075 85.090 203.135 ;
        RECT 84.770 202.935 85.920 203.075 ;
        RECT 84.770 202.875 85.090 202.935 ;
        RECT 79.710 202.735 80.030 202.795 ;
        RECT 80.185 202.735 80.475 202.780 ;
        RECT 79.710 202.595 80.475 202.735 ;
        RECT 79.710 202.535 80.030 202.595 ;
        RECT 80.185 202.550 80.475 202.595 ;
        RECT 83.390 202.535 83.710 202.795 ;
        RECT 84.325 202.735 84.615 202.780 ;
        RECT 85.230 202.735 85.550 202.795 ;
        RECT 85.780 202.780 85.920 202.935 ;
        RECT 87.070 202.875 87.390 203.135 ;
        RECT 88.540 202.780 88.680 203.615 ;
        RECT 106.850 203.555 107.170 203.615 ;
        RECT 107.310 203.755 107.630 203.815 ;
        RECT 109.150 203.755 109.470 203.815 ;
        RECT 116.970 203.755 117.290 203.815 ;
        RECT 107.310 203.615 117.290 203.755 ;
        RECT 107.310 203.555 107.630 203.615 ;
        RECT 109.150 203.555 109.470 203.615 ;
        RECT 88.910 203.415 89.230 203.475 ;
        RECT 96.730 203.415 97.050 203.475 ;
        RECT 99.490 203.415 99.810 203.475 ;
        RECT 104.090 203.415 104.410 203.475 ;
        RECT 110.085 203.415 110.375 203.460 ;
        RECT 88.910 203.275 91.440 203.415 ;
        RECT 88.910 203.215 89.230 203.275 ;
        RECT 84.325 202.595 85.550 202.735 ;
        RECT 84.325 202.550 84.615 202.595 ;
        RECT 85.230 202.535 85.550 202.595 ;
        RECT 85.705 202.550 85.995 202.780 ;
        RECT 88.465 202.550 88.755 202.780 ;
        RECT 88.910 202.535 89.230 202.795 ;
        RECT 89.370 202.735 89.690 202.795 ;
        RECT 91.300 202.780 91.440 203.275 ;
        RECT 95.900 203.275 97.050 203.415 ;
        RECT 93.970 203.075 94.290 203.135 ;
        RECT 92.220 202.935 94.290 203.075 ;
        RECT 89.845 202.735 90.135 202.780 ;
        RECT 89.370 202.595 90.135 202.735 ;
        RECT 89.370 202.535 89.690 202.595 ;
        RECT 89.845 202.550 90.135 202.595 ;
        RECT 90.305 202.550 90.595 202.780 ;
        RECT 91.225 202.735 91.515 202.780 ;
        RECT 91.670 202.735 91.990 202.795 ;
        RECT 92.220 202.780 92.360 202.935 ;
        RECT 93.970 202.875 94.290 202.935 ;
        RECT 91.225 202.595 91.990 202.735 ;
        RECT 91.225 202.550 91.515 202.595 ;
        RECT 90.380 202.395 90.520 202.550 ;
        RECT 91.670 202.535 91.990 202.595 ;
        RECT 92.145 202.550 92.435 202.780 ;
        RECT 93.065 202.550 93.355 202.780 ;
        RECT 79.340 202.255 90.520 202.395 ;
        RECT 93.140 202.395 93.280 202.550 ;
        RECT 93.510 202.535 93.830 202.795 ;
        RECT 95.900 202.780 96.040 203.275 ;
        RECT 96.730 203.215 97.050 203.275 ;
        RECT 97.280 203.275 99.810 203.415 ;
        RECT 97.280 203.075 97.420 203.275 ;
        RECT 99.490 203.215 99.810 203.275 ;
        RECT 100.960 203.275 103.400 203.415 ;
        RECT 100.960 203.075 101.100 203.275 ;
        RECT 96.360 202.935 97.420 203.075 ;
        RECT 97.740 202.935 101.100 203.075 ;
        RECT 96.360 202.795 96.500 202.935 ;
        RECT 97.740 202.795 97.880 202.935 ;
        RECT 94.445 202.735 94.735 202.780 ;
        RECT 94.905 202.735 95.195 202.780 ;
        RECT 94.445 202.595 95.195 202.735 ;
        RECT 94.445 202.550 94.735 202.595 ;
        RECT 94.905 202.550 95.195 202.595 ;
        RECT 95.825 202.550 96.115 202.780 ;
        RECT 96.270 202.535 96.590 202.795 ;
        RECT 97.190 202.535 97.510 202.795 ;
        RECT 97.650 202.535 97.970 202.795 ;
        RECT 98.570 202.735 98.890 202.795 ;
        RECT 99.045 202.735 99.335 202.780 ;
        RECT 98.570 202.595 99.335 202.735 ;
        RECT 98.570 202.535 98.890 202.595 ;
        RECT 99.045 202.550 99.335 202.595 ;
        RECT 98.125 202.395 98.415 202.440 ;
        RECT 93.140 202.255 98.415 202.395 ;
        RECT 99.120 202.395 99.260 202.550 ;
        RECT 99.490 202.535 99.810 202.795 ;
        RECT 100.410 202.535 100.730 202.795 ;
        RECT 100.960 202.780 101.100 202.935 ;
        RECT 101.330 203.075 101.650 203.135 ;
        RECT 103.260 203.075 103.400 203.275 ;
        RECT 104.090 203.275 110.375 203.415 ;
        RECT 104.090 203.215 104.410 203.275 ;
        RECT 110.085 203.230 110.375 203.275 ;
        RECT 107.325 203.075 107.615 203.120 ;
        RECT 101.330 202.935 102.940 203.075 ;
        RECT 103.260 202.935 107.615 203.075 ;
        RECT 101.330 202.875 101.650 202.935 ;
        RECT 100.885 202.550 101.175 202.780 ;
        RECT 102.250 202.535 102.570 202.795 ;
        RECT 102.800 202.735 102.940 202.935 ;
        RECT 107.325 202.890 107.615 202.935 ;
        RECT 107.770 203.075 108.090 203.135 ;
        RECT 111.450 203.075 111.770 203.135 ;
        RECT 112.000 203.120 112.140 203.615 ;
        RECT 116.970 203.555 117.290 203.615 ;
        RECT 118.350 203.555 118.670 203.815 ;
        RECT 120.740 203.615 142.960 203.755 ;
        RECT 113.750 203.215 114.070 203.475 ;
        RECT 117.445 203.415 117.735 203.460 ;
        RECT 120.740 203.415 120.880 203.615 ;
        RECT 117.445 203.275 120.880 203.415 ;
        RECT 121.225 203.415 121.515 203.460 ;
        RECT 124.345 203.415 124.635 203.460 ;
        RECT 126.235 203.415 126.525 203.460 ;
        RECT 121.225 203.275 126.525 203.415 ;
        RECT 117.445 203.230 117.735 203.275 ;
        RECT 121.225 203.230 121.515 203.275 ;
        RECT 124.345 203.230 124.635 203.275 ;
        RECT 126.235 203.230 126.525 203.275 ;
        RECT 128.470 203.415 128.790 203.475 ;
        RECT 130.325 203.415 130.615 203.460 ;
        RECT 128.470 203.275 130.615 203.415 ;
        RECT 128.470 203.215 128.790 203.275 ;
        RECT 130.325 203.230 130.615 203.275 ;
        RECT 133.185 203.415 133.475 203.460 ;
        RECT 136.305 203.415 136.595 203.460 ;
        RECT 138.195 203.415 138.485 203.460 ;
        RECT 133.185 203.275 138.485 203.415 ;
        RECT 133.185 203.230 133.475 203.275 ;
        RECT 136.305 203.230 136.595 203.275 ;
        RECT 138.195 203.230 138.485 203.275 ;
        RECT 107.770 202.935 111.770 203.075 ;
        RECT 107.770 202.875 108.090 202.935 ;
        RECT 111.450 202.875 111.770 202.935 ;
        RECT 111.925 202.890 112.215 203.120 ;
        RECT 112.385 203.075 112.675 203.120 ;
        RECT 122.030 203.075 122.350 203.135 ;
        RECT 127.105 203.075 127.395 203.120 ;
        RECT 112.385 202.935 115.820 203.075 ;
        RECT 112.385 202.890 112.675 202.935 ;
        RECT 103.185 202.735 103.475 202.780 ;
        RECT 102.800 202.595 103.475 202.735 ;
        RECT 103.185 202.550 103.475 202.595 ;
        RECT 104.550 202.535 104.870 202.795 ;
        RECT 106.850 202.535 107.170 202.795 ;
        RECT 109.610 202.535 109.930 202.795 ;
        RECT 110.070 202.735 110.390 202.795 ;
        RECT 111.005 202.735 111.295 202.780 ;
        RECT 112.830 202.735 113.150 202.795 ;
        RECT 110.070 202.595 113.150 202.735 ;
        RECT 110.070 202.535 110.390 202.595 ;
        RECT 111.005 202.550 111.295 202.595 ;
        RECT 112.830 202.535 113.150 202.595 ;
        RECT 113.305 202.550 113.595 202.780 ;
        RECT 104.640 202.395 104.780 202.535 ;
        RECT 106.405 202.395 106.695 202.440 ;
        RECT 109.165 202.395 109.455 202.440 ;
        RECT 99.120 202.255 109.455 202.395 ;
        RECT 25.890 202.055 26.210 202.115 ;
        RECT 26.810 202.055 27.130 202.115 ;
        RECT 29.585 202.055 29.875 202.100 ;
        RECT 25.890 201.915 29.875 202.055 ;
        RECT 25.890 201.855 26.210 201.915 ;
        RECT 26.810 201.855 27.130 201.915 ;
        RECT 29.585 201.870 29.875 201.915 ;
        RECT 32.790 202.055 33.110 202.115 ;
        RECT 38.310 202.055 38.630 202.115 ;
        RECT 32.790 201.915 38.630 202.055 ;
        RECT 32.790 201.855 33.110 201.915 ;
        RECT 38.310 201.855 38.630 201.915 ;
        RECT 43.830 201.855 44.150 202.115 ;
        RECT 44.750 202.055 45.070 202.115 ;
        RECT 54.040 202.055 54.180 202.210 ;
        RECT 44.750 201.915 54.180 202.055 ;
        RECT 55.420 202.055 55.560 202.210 ;
        RECT 69.130 202.195 69.450 202.255 ;
        RECT 98.125 202.210 98.415 202.255 ;
        RECT 106.405 202.210 106.695 202.255 ;
        RECT 109.165 202.210 109.455 202.255 ;
        RECT 57.170 202.055 57.490 202.115 ;
        RECT 55.420 201.915 57.490 202.055 ;
        RECT 44.750 201.855 45.070 201.915 ;
        RECT 57.170 201.855 57.490 201.915 ;
        RECT 60.405 202.055 60.695 202.100 ;
        RECT 62.690 202.055 63.010 202.115 ;
        RECT 60.405 201.915 63.010 202.055 ;
        RECT 60.405 201.870 60.695 201.915 ;
        RECT 62.690 201.855 63.010 201.915 ;
        RECT 68.210 202.055 68.530 202.115 ;
        RECT 70.065 202.055 70.355 202.100 ;
        RECT 68.210 201.915 70.355 202.055 ;
        RECT 68.210 201.855 68.530 201.915 ;
        RECT 70.065 201.870 70.355 201.915 ;
        RECT 76.965 202.055 77.255 202.100 ;
        RECT 82.470 202.055 82.790 202.115 ;
        RECT 76.965 201.915 82.790 202.055 ;
        RECT 76.965 201.870 77.255 201.915 ;
        RECT 82.470 201.855 82.790 201.915 ;
        RECT 84.770 202.055 85.090 202.115 ;
        RECT 88.910 202.055 89.230 202.115 ;
        RECT 84.770 201.915 89.230 202.055 ;
        RECT 84.770 201.855 85.090 201.915 ;
        RECT 88.910 201.855 89.230 201.915 ;
        RECT 89.370 201.855 89.690 202.115 ;
        RECT 90.750 201.855 91.070 202.115 ;
        RECT 92.130 201.855 92.450 202.115 ;
        RECT 93.510 201.855 93.830 202.115 ;
        RECT 97.190 202.055 97.510 202.115 ;
        RECT 100.410 202.055 100.730 202.115 ;
        RECT 97.190 201.915 100.730 202.055 ;
        RECT 97.190 201.855 97.510 201.915 ;
        RECT 100.410 201.855 100.730 201.915 ;
        RECT 101.330 202.055 101.650 202.115 ;
        RECT 102.710 202.055 103.030 202.115 ;
        RECT 101.330 201.915 103.030 202.055 ;
        RECT 101.330 201.855 101.650 201.915 ;
        RECT 102.710 201.855 103.030 201.915 ;
        RECT 103.185 202.055 103.475 202.100 ;
        RECT 103.630 202.055 103.950 202.115 ;
        RECT 103.185 201.915 103.950 202.055 ;
        RECT 103.185 201.870 103.475 201.915 ;
        RECT 103.630 201.855 103.950 201.915 ;
        RECT 104.090 202.055 104.410 202.115 ;
        RECT 104.565 202.055 104.855 202.100 ;
        RECT 104.090 201.915 104.855 202.055 ;
        RECT 104.090 201.855 104.410 201.915 ;
        RECT 104.565 201.870 104.855 201.915 ;
        RECT 105.470 202.055 105.790 202.115 ;
        RECT 113.380 202.055 113.520 202.550 ;
        RECT 114.210 202.535 114.530 202.795 ;
        RECT 114.670 202.535 114.990 202.795 ;
        RECT 105.470 201.915 113.520 202.055 ;
        RECT 114.760 202.055 114.900 202.535 ;
        RECT 115.680 202.455 115.820 202.935 ;
        RECT 122.030 202.935 139.280 203.075 ;
        RECT 122.030 202.875 122.350 202.935 ;
        RECT 127.105 202.890 127.395 202.935 ;
        RECT 116.510 202.535 116.830 202.795 ;
        RECT 115.590 202.195 115.910 202.455 ;
        RECT 116.065 202.395 116.355 202.440 ;
        RECT 116.970 202.395 117.290 202.455 ;
        RECT 118.810 202.395 119.130 202.455 ;
        RECT 120.145 202.440 120.435 202.755 ;
        RECT 121.225 202.735 121.515 202.780 ;
        RECT 124.805 202.735 125.095 202.780 ;
        RECT 126.640 202.735 126.930 202.780 ;
        RECT 121.225 202.595 126.930 202.735 ;
        RECT 121.225 202.550 121.515 202.595 ;
        RECT 124.805 202.550 125.095 202.595 ;
        RECT 126.640 202.550 126.930 202.595 ;
        RECT 128.470 202.535 128.790 202.795 ;
        RECT 129.405 202.735 129.695 202.780 ;
        RECT 129.850 202.735 130.170 202.795 ;
        RECT 139.140 202.780 139.280 202.935 ;
        RECT 142.820 202.780 142.960 203.615 ;
        RECT 145.490 203.555 145.810 203.815 ;
        RECT 129.405 202.595 130.170 202.735 ;
        RECT 129.405 202.550 129.695 202.595 ;
        RECT 129.850 202.535 130.170 202.595 ;
        RECT 116.065 202.255 119.130 202.395 ;
        RECT 116.065 202.210 116.355 202.255 ;
        RECT 116.970 202.195 117.290 202.255 ;
        RECT 118.810 202.195 119.130 202.255 ;
        RECT 119.845 202.395 120.435 202.440 ;
        RECT 123.085 202.395 123.735 202.440 ;
        RECT 119.845 202.255 125.015 202.395 ;
        RECT 119.845 202.210 120.135 202.255 ;
        RECT 123.085 202.210 123.735 202.255 ;
        RECT 124.330 202.055 124.650 202.115 ;
        RECT 114.760 201.915 124.650 202.055 ;
        RECT 124.875 202.055 125.015 202.255 ;
        RECT 125.710 202.195 126.030 202.455 ;
        RECT 132.105 202.440 132.395 202.755 ;
        RECT 133.185 202.735 133.475 202.780 ;
        RECT 136.765 202.735 137.055 202.780 ;
        RECT 138.600 202.735 138.890 202.780 ;
        RECT 133.185 202.595 138.890 202.735 ;
        RECT 133.185 202.550 133.475 202.595 ;
        RECT 136.765 202.550 137.055 202.595 ;
        RECT 138.600 202.550 138.890 202.595 ;
        RECT 139.065 202.735 139.355 202.780 ;
        RECT 139.525 202.735 139.815 202.780 ;
        RECT 139.065 202.595 139.815 202.735 ;
        RECT 139.065 202.550 139.355 202.595 ;
        RECT 139.525 202.550 139.815 202.595 ;
        RECT 141.365 202.550 141.655 202.780 ;
        RECT 142.745 202.550 143.035 202.780 ;
        RECT 144.585 202.735 144.875 202.780 ;
        RECT 145.030 202.735 145.350 202.795 ;
        RECT 144.585 202.595 145.350 202.735 ;
        RECT 144.585 202.550 144.875 202.595 ;
        RECT 131.805 202.395 132.395 202.440 ;
        RECT 133.990 202.395 134.310 202.455 ;
        RECT 135.045 202.395 135.695 202.440 ;
        RECT 131.805 202.255 135.695 202.395 ;
        RECT 131.805 202.210 132.095 202.255 ;
        RECT 133.990 202.195 134.310 202.255 ;
        RECT 135.045 202.210 135.695 202.255 ;
        RECT 137.685 202.210 137.975 202.440 ;
        RECT 141.440 202.395 141.580 202.550 ;
        RECT 145.030 202.535 145.350 202.595 ;
        RECT 138.680 202.255 141.580 202.395 ;
        RECT 126.630 202.055 126.950 202.115 ;
        RECT 124.875 201.915 126.950 202.055 ;
        RECT 105.470 201.855 105.790 201.915 ;
        RECT 124.330 201.855 124.650 201.915 ;
        RECT 126.630 201.855 126.950 201.915 ;
        RECT 127.565 202.055 127.855 202.100 ;
        RECT 129.390 202.055 129.710 202.115 ;
        RECT 127.565 201.915 129.710 202.055 ;
        RECT 127.565 201.870 127.855 201.915 ;
        RECT 129.390 201.855 129.710 201.915 ;
        RECT 130.770 202.055 131.090 202.115 ;
        RECT 137.760 202.055 137.900 202.210 ;
        RECT 138.680 202.115 138.820 202.255 ;
        RECT 130.770 201.915 137.900 202.055 ;
        RECT 130.770 201.855 131.090 201.915 ;
        RECT 138.590 201.855 138.910 202.115 ;
        RECT 139.970 201.855 140.290 202.115 ;
        RECT 142.285 202.055 142.575 202.100 ;
        RECT 143.190 202.055 143.510 202.115 ;
        RECT 142.285 201.915 143.510 202.055 ;
        RECT 142.285 201.870 142.575 201.915 ;
        RECT 143.190 201.855 143.510 201.915 ;
        RECT 143.650 201.855 143.970 202.115 ;
        RECT 13.860 201.235 147.720 201.715 ;
        RECT 28.650 201.035 28.970 201.095 ;
        RECT 36.930 201.035 37.250 201.095 ;
        RECT 28.650 200.895 37.250 201.035 ;
        RECT 28.650 200.835 28.970 200.895 ;
        RECT 36.930 200.835 37.250 200.895 ;
        RECT 40.150 200.835 40.470 201.095 ;
        RECT 43.845 201.035 44.135 201.080 ;
        RECT 45.670 201.035 45.990 201.095 ;
        RECT 43.845 200.895 45.990 201.035 ;
        RECT 43.845 200.850 44.135 200.895 ;
        RECT 45.670 200.835 45.990 200.895 ;
        RECT 48.430 201.035 48.750 201.095 ;
        RECT 61.310 201.035 61.630 201.095 ;
        RECT 63.625 201.035 63.915 201.080 ;
        RECT 64.990 201.035 65.310 201.095 ;
        RECT 48.430 200.895 61.630 201.035 ;
        RECT 48.430 200.835 48.750 200.895 ;
        RECT 61.310 200.835 61.630 200.895 ;
        RECT 62.320 200.895 65.310 201.035 ;
        RECT 23.125 200.695 23.775 200.740 ;
        RECT 26.725 200.695 27.015 200.740 ;
        RECT 23.125 200.555 27.015 200.695 ;
        RECT 23.125 200.510 23.775 200.555 ;
        RECT 26.425 200.510 27.015 200.555 ;
        RECT 32.805 200.695 33.095 200.740 ;
        RECT 33.250 200.695 33.570 200.755 ;
        RECT 34.630 200.695 34.950 200.755 ;
        RECT 44.765 200.695 45.055 200.740 ;
        RECT 45.210 200.695 45.530 200.755 ;
        RECT 53.490 200.695 53.810 200.755 ;
        RECT 32.805 200.555 34.950 200.695 ;
        RECT 32.805 200.510 33.095 200.555 ;
        RECT 26.425 200.415 26.715 200.510 ;
        RECT 33.250 200.495 33.570 200.555 ;
        RECT 34.630 200.495 34.950 200.555 ;
        RECT 37.940 200.555 44.060 200.695 ;
        RECT 16.705 200.355 16.995 200.400 ;
        RECT 18.070 200.355 18.390 200.415 ;
        RECT 16.705 200.215 18.390 200.355 ;
        RECT 16.705 200.170 16.995 200.215 ;
        RECT 18.070 200.155 18.390 200.215 ;
        RECT 18.545 200.170 18.835 200.400 ;
        RECT 18.990 200.355 19.310 200.415 ;
        RECT 19.465 200.355 19.755 200.400 ;
        RECT 18.990 200.215 19.755 200.355 ;
        RECT 15.770 199.475 16.090 199.735 ;
        RECT 17.610 199.475 17.930 199.735 ;
        RECT 18.620 199.675 18.760 200.170 ;
        RECT 18.990 200.155 19.310 200.215 ;
        RECT 19.465 200.170 19.755 200.215 ;
        RECT 19.930 200.355 20.220 200.400 ;
        RECT 21.765 200.355 22.055 200.400 ;
        RECT 25.345 200.355 25.635 200.400 ;
        RECT 19.930 200.215 25.635 200.355 ;
        RECT 19.930 200.170 20.220 200.215 ;
        RECT 21.765 200.170 22.055 200.215 ;
        RECT 25.345 200.170 25.635 200.215 ;
        RECT 26.350 200.195 26.715 200.415 ;
        RECT 30.030 200.355 30.350 200.415 ;
        RECT 30.505 200.355 30.795 200.400 ;
        RECT 30.950 200.355 31.270 200.415 ;
        RECT 30.030 200.215 31.270 200.355 ;
        RECT 26.350 200.155 26.670 200.195 ;
        RECT 30.030 200.155 30.350 200.215 ;
        RECT 30.505 200.170 30.795 200.215 ;
        RECT 30.950 200.155 31.270 200.215 ;
        RECT 31.410 200.155 31.730 200.415 ;
        RECT 33.725 200.355 34.015 200.400 ;
        RECT 34.170 200.355 34.490 200.415 ;
        RECT 33.725 200.215 34.490 200.355 ;
        RECT 33.725 200.170 34.015 200.215 ;
        RECT 34.170 200.155 34.490 200.215 ;
        RECT 35.550 200.400 35.870 200.415 ;
        RECT 35.550 200.170 36.085 200.400 ;
        RECT 35.550 200.155 35.870 200.170 ;
        RECT 36.470 200.155 36.790 200.415 ;
        RECT 36.930 200.155 37.250 200.415 ;
        RECT 37.390 200.355 37.710 200.415 ;
        RECT 37.940 200.400 38.080 200.555 ;
        RECT 41.070 200.400 41.390 200.415 ;
        RECT 37.860 200.355 38.150 200.400 ;
        RECT 37.390 200.215 38.150 200.355 ;
        RECT 37.390 200.155 37.710 200.215 ;
        RECT 37.860 200.170 38.150 200.215 ;
        RECT 38.325 200.170 38.615 200.400 ;
        RECT 41.060 200.355 41.390 200.400 ;
        RECT 40.875 200.215 41.390 200.355 ;
        RECT 41.060 200.170 41.390 200.215 ;
        RECT 20.845 200.015 21.135 200.060 ;
        RECT 27.270 200.015 27.590 200.075 ;
        RECT 20.845 199.875 27.590 200.015 ;
        RECT 20.845 199.830 21.135 199.875 ;
        RECT 27.270 199.815 27.590 199.875 ;
        RECT 28.190 200.015 28.510 200.075 ;
        RECT 29.585 200.015 29.875 200.060 ;
        RECT 28.190 199.875 29.875 200.015 ;
        RECT 28.190 199.815 28.510 199.875 ;
        RECT 29.585 199.830 29.875 199.875 ;
        RECT 32.345 200.015 32.635 200.060 ;
        RECT 38.400 200.015 38.540 200.170 ;
        RECT 41.070 200.155 41.390 200.170 ;
        RECT 41.530 200.155 41.850 200.415 ;
        RECT 42.005 200.170 42.295 200.400 ;
        RECT 42.450 200.355 42.770 200.415 ;
        RECT 42.920 200.355 43.210 200.400 ;
        RECT 42.450 200.215 43.210 200.355 ;
        RECT 32.345 199.875 38.540 200.015 ;
        RECT 42.080 200.015 42.220 200.170 ;
        RECT 42.450 200.155 42.770 200.215 ;
        RECT 42.920 200.170 43.210 200.215 ;
        RECT 43.385 200.170 43.675 200.400 ;
        RECT 43.920 200.355 44.060 200.555 ;
        RECT 44.765 200.555 46.360 200.695 ;
        RECT 44.765 200.510 45.055 200.555 ;
        RECT 45.210 200.495 45.530 200.555 ;
        RECT 45.670 200.355 45.990 200.415 ;
        RECT 46.220 200.400 46.360 200.555 ;
        RECT 48.980 200.555 53.810 200.695 ;
        RECT 43.920 200.215 45.990 200.355 ;
        RECT 43.460 200.015 43.600 200.170 ;
        RECT 45.670 200.155 45.990 200.215 ;
        RECT 46.145 200.170 46.435 200.400 ;
        RECT 47.065 200.170 47.355 200.400 ;
        RECT 46.605 200.015 46.895 200.060 ;
        RECT 42.080 199.875 43.140 200.015 ;
        RECT 43.460 199.875 46.895 200.015 ;
        RECT 32.345 199.830 32.635 199.875 ;
        RECT 19.450 199.675 19.770 199.735 ;
        RECT 18.620 199.535 19.770 199.675 ;
        RECT 19.450 199.475 19.770 199.535 ;
        RECT 20.335 199.675 20.625 199.720 ;
        RECT 22.225 199.675 22.515 199.720 ;
        RECT 25.345 199.675 25.635 199.720 ;
        RECT 20.335 199.535 25.635 199.675 ;
        RECT 20.335 199.490 20.625 199.535 ;
        RECT 22.225 199.490 22.515 199.535 ;
        RECT 25.345 199.490 25.635 199.535 ;
        RECT 34.645 199.675 34.935 199.720 ;
        RECT 42.450 199.675 42.770 199.735 ;
        RECT 34.645 199.535 42.770 199.675 ;
        RECT 43.000 199.675 43.140 199.875 ;
        RECT 46.605 199.830 46.895 199.875 ;
        RECT 43.370 199.675 43.690 199.735 ;
        RECT 43.000 199.535 43.690 199.675 ;
        RECT 34.645 199.490 34.935 199.535 ;
        RECT 42.450 199.475 42.770 199.535 ;
        RECT 43.370 199.475 43.690 199.535 ;
        RECT 43.830 199.675 44.150 199.735 ;
        RECT 47.140 199.675 47.280 200.170 ;
        RECT 48.430 200.155 48.750 200.415 ;
        RECT 48.980 200.400 49.120 200.555 ;
        RECT 50.820 200.400 50.960 200.555 ;
        RECT 53.490 200.495 53.810 200.555 ;
        RECT 55.805 200.695 56.095 200.740 ;
        RECT 57.630 200.695 57.950 200.755 ;
        RECT 61.770 200.695 62.090 200.755 ;
        RECT 55.805 200.555 57.950 200.695 ;
        RECT 55.805 200.510 56.095 200.555 ;
        RECT 57.630 200.495 57.950 200.555 ;
        RECT 59.560 200.555 62.090 200.695 ;
        RECT 48.905 200.170 49.195 200.400 ;
        RECT 49.825 200.355 50.115 200.400 ;
        RECT 49.440 200.215 50.115 200.355 ;
        RECT 47.510 199.815 47.830 200.075 ;
        RECT 49.440 200.015 49.580 200.215 ;
        RECT 49.825 200.170 50.115 200.215 ;
        RECT 50.285 200.170 50.575 200.400 ;
        RECT 50.745 200.170 51.035 200.400 ;
        RECT 52.125 200.170 52.415 200.400 ;
        RECT 54.425 200.170 54.715 200.400 ;
        RECT 54.885 200.170 55.175 200.400 ;
        RECT 48.980 199.875 49.580 200.015 ;
        RECT 50.360 200.015 50.500 200.170 ;
        RECT 51.650 200.015 51.970 200.075 ;
        RECT 52.200 200.015 52.340 200.170 ;
        RECT 50.360 199.875 50.960 200.015 ;
        RECT 43.830 199.535 47.280 199.675 ;
        RECT 48.980 199.675 49.120 199.875 ;
        RECT 50.270 199.675 50.590 199.735 ;
        RECT 48.980 199.535 50.590 199.675 ;
        RECT 43.830 199.475 44.150 199.535 ;
        RECT 24.050 199.335 24.370 199.395 ;
        RECT 35.105 199.335 35.395 199.380 ;
        RECT 24.050 199.195 35.395 199.335 ;
        RECT 24.050 199.135 24.370 199.195 ;
        RECT 35.105 199.150 35.395 199.195 ;
        RECT 36.470 199.335 36.790 199.395 ;
        RECT 41.530 199.335 41.850 199.395 ;
        RECT 43.920 199.335 44.060 199.475 ;
        RECT 36.470 199.195 44.060 199.335 ;
        RECT 47.140 199.335 47.280 199.535 ;
        RECT 50.270 199.475 50.590 199.535 ;
        RECT 50.820 199.675 50.960 199.875 ;
        RECT 51.650 199.875 52.340 200.015 ;
        RECT 51.650 199.815 51.970 199.875 ;
        RECT 52.570 199.815 52.890 200.075 ;
        RECT 54.500 199.675 54.640 200.170 ;
        RECT 54.960 200.015 55.100 200.170 ;
        RECT 55.330 200.155 55.650 200.415 ;
        RECT 56.710 200.155 57.030 200.415 ;
        RECT 59.560 200.400 59.700 200.555 ;
        RECT 61.770 200.495 62.090 200.555 ;
        RECT 58.105 200.355 58.395 200.400 ;
        RECT 57.260 200.215 58.395 200.355 ;
        RECT 57.260 200.015 57.400 200.215 ;
        RECT 58.105 200.170 58.395 200.215 ;
        RECT 58.570 200.170 58.860 200.400 ;
        RECT 59.485 200.170 59.775 200.400 ;
        RECT 54.960 199.875 57.400 200.015 ;
        RECT 57.645 200.015 57.935 200.060 ;
        RECT 58.640 200.015 58.780 200.170 ;
        RECT 59.930 200.155 60.250 200.415 ;
        RECT 60.635 200.355 60.925 200.400 ;
        RECT 62.320 200.355 62.460 200.895 ;
        RECT 63.625 200.850 63.915 200.895 ;
        RECT 64.990 200.835 65.310 200.895 ;
        RECT 65.925 201.035 66.215 201.080 ;
        RECT 68.670 201.035 68.990 201.095 ;
        RECT 65.925 200.895 68.990 201.035 ;
        RECT 65.925 200.850 66.215 200.895 ;
        RECT 68.670 200.835 68.990 200.895 ;
        RECT 69.130 201.035 69.450 201.095 ;
        RECT 70.970 201.035 71.290 201.095 ;
        RECT 69.130 200.895 71.290 201.035 ;
        RECT 69.130 200.835 69.450 200.895 ;
        RECT 70.970 200.835 71.290 200.895 ;
        RECT 73.285 201.035 73.575 201.080 ;
        RECT 76.030 201.035 76.350 201.095 ;
        RECT 97.650 201.035 97.970 201.095 ;
        RECT 73.285 200.895 76.350 201.035 ;
        RECT 73.285 200.850 73.575 200.895 ;
        RECT 76.030 200.835 76.350 200.895 ;
        RECT 79.800 200.895 97.970 201.035 ;
        RECT 79.800 200.755 79.940 200.895 ;
        RECT 97.650 200.835 97.970 200.895 ;
        RECT 98.110 201.035 98.430 201.095 ;
        RECT 99.490 201.035 99.810 201.095 ;
        RECT 105.010 201.035 105.330 201.095 ;
        RECT 109.150 201.035 109.470 201.095 ;
        RECT 122.030 201.035 122.350 201.095 ;
        RECT 98.110 200.895 98.800 201.035 ;
        RECT 98.110 200.835 98.430 200.895 ;
        RECT 73.730 200.695 74.050 200.755 ;
        RECT 70.600 200.555 74.050 200.695 ;
        RECT 70.600 200.415 70.740 200.555 ;
        RECT 73.730 200.495 74.050 200.555 ;
        RECT 74.665 200.695 74.955 200.740 ;
        RECT 76.490 200.695 76.810 200.755 ;
        RECT 79.710 200.695 80.030 200.755 ;
        RECT 83.390 200.695 83.710 200.755 ;
        RECT 74.665 200.555 76.810 200.695 ;
        RECT 74.665 200.510 74.955 200.555 ;
        RECT 76.490 200.495 76.810 200.555 ;
        RECT 77.500 200.555 80.030 200.695 ;
        RECT 60.635 200.215 62.460 200.355 ;
        RECT 60.635 200.170 60.925 200.215 ;
        RECT 62.690 200.155 63.010 200.415 ;
        RECT 64.070 200.155 64.390 200.415 ;
        RECT 66.845 200.355 67.135 200.400 ;
        RECT 67.290 200.355 67.610 200.415 ;
        RECT 66.845 200.215 67.610 200.355 ;
        RECT 66.845 200.170 67.135 200.215 ;
        RECT 67.290 200.155 67.610 200.215 ;
        RECT 67.765 200.170 68.055 200.400 ;
        RECT 57.645 199.875 58.780 200.015 ;
        RECT 57.645 199.830 57.935 199.875 ;
        RECT 61.770 199.815 62.090 200.075 ;
        RECT 63.610 200.015 63.930 200.075 ;
        RECT 66.370 200.015 66.690 200.075 ;
        RECT 63.610 199.875 66.690 200.015 ;
        RECT 67.840 200.015 67.980 200.170 ;
        RECT 68.210 200.155 68.530 200.415 ;
        RECT 69.590 200.155 69.910 200.415 ;
        RECT 70.065 200.170 70.355 200.400 ;
        RECT 68.685 200.015 68.975 200.060 ;
        RECT 67.840 199.875 68.975 200.015 ;
        RECT 70.140 200.015 70.280 200.170 ;
        RECT 70.510 200.155 70.830 200.415 ;
        RECT 70.970 200.355 71.290 200.415 ;
        RECT 71.445 200.355 71.735 200.400 ;
        RECT 70.970 200.215 71.735 200.355 ;
        RECT 70.970 200.155 71.290 200.215 ;
        RECT 71.445 200.170 71.735 200.215 ;
        RECT 72.350 200.155 72.670 200.415 ;
        RECT 75.585 200.355 75.875 200.400 ;
        RECT 74.740 200.215 75.875 200.355 ;
        RECT 72.440 200.015 72.580 200.155 ;
        RECT 74.740 200.075 74.880 200.215 ;
        RECT 75.585 200.170 75.875 200.215 ;
        RECT 76.045 200.355 76.335 200.400 ;
        RECT 76.045 200.215 76.720 200.355 ;
        RECT 76.045 200.170 76.335 200.215 ;
        RECT 70.140 199.875 72.580 200.015 ;
        RECT 63.610 199.815 63.930 199.875 ;
        RECT 66.370 199.815 66.690 199.875 ;
        RECT 68.685 199.830 68.975 199.875 ;
        RECT 74.650 199.815 74.970 200.075 ;
        RECT 76.580 200.015 76.720 200.215 ;
        RECT 76.950 200.155 77.270 200.415 ;
        RECT 77.500 200.400 77.640 200.555 ;
        RECT 79.710 200.495 80.030 200.555 ;
        RECT 80.260 200.555 83.710 200.695 ;
        RECT 77.425 200.170 77.715 200.400 ;
        RECT 78.790 200.155 79.110 200.415 ;
        RECT 80.260 200.400 80.400 200.555 ;
        RECT 83.390 200.495 83.710 200.555 ;
        RECT 84.310 200.695 84.630 200.755 ;
        RECT 90.290 200.695 90.610 200.755 ;
        RECT 93.065 200.695 93.355 200.740 ;
        RECT 95.810 200.695 96.130 200.755 ;
        RECT 98.660 200.740 98.800 200.895 ;
        RECT 99.490 200.895 105.330 201.035 ;
        RECT 99.490 200.835 99.810 200.895 ;
        RECT 105.010 200.835 105.330 200.895 ;
        RECT 107.400 200.895 109.470 201.035 ;
        RECT 84.310 200.555 96.130 200.695 ;
        RECT 84.310 200.495 84.630 200.555 ;
        RECT 80.185 200.170 80.475 200.400 ;
        RECT 81.090 200.355 81.410 200.415 ;
        RECT 82.485 200.355 82.775 200.400 ;
        RECT 81.090 200.215 82.775 200.355 ;
        RECT 81.090 200.155 81.410 200.215 ;
        RECT 82.485 200.170 82.775 200.215 ;
        RECT 84.785 200.170 85.075 200.400 ;
        RECT 76.580 199.875 77.640 200.015 ;
        RECT 56.710 199.675 57.030 199.735 ;
        RECT 50.820 199.535 57.030 199.675 ;
        RECT 47.970 199.335 48.290 199.395 ;
        RECT 50.820 199.335 50.960 199.535 ;
        RECT 56.710 199.475 57.030 199.535 ;
        RECT 58.090 199.675 58.410 199.735 ;
        RECT 61.325 199.675 61.615 199.720 ;
        RECT 58.090 199.535 61.615 199.675 ;
        RECT 58.090 199.475 58.410 199.535 ;
        RECT 61.325 199.490 61.615 199.535 ;
        RECT 62.230 199.675 62.550 199.735 ;
        RECT 74.740 199.675 74.880 199.815 ;
        RECT 77.500 199.675 77.640 199.875 ;
        RECT 77.870 199.815 78.190 200.075 ;
        RECT 79.265 199.830 79.555 200.060 ;
        RECT 79.340 199.675 79.480 199.830 ;
        RECT 79.710 199.815 80.030 200.075 ;
        RECT 80.630 200.015 80.950 200.075 ;
        RECT 81.565 200.015 81.855 200.060 ;
        RECT 80.630 199.875 81.855 200.015 ;
        RECT 80.630 199.815 80.950 199.875 ;
        RECT 81.565 199.830 81.855 199.875 ;
        RECT 83.405 199.830 83.695 200.060 ;
        RECT 62.230 199.535 73.500 199.675 ;
        RECT 74.740 199.535 77.180 199.675 ;
        RECT 77.500 199.535 80.400 199.675 ;
        RECT 62.230 199.475 62.550 199.535 ;
        RECT 47.140 199.195 50.960 199.335 ;
        RECT 51.205 199.335 51.495 199.380 ;
        RECT 56.250 199.335 56.570 199.395 ;
        RECT 71.445 199.335 71.735 199.380 ;
        RECT 51.205 199.195 71.735 199.335 ;
        RECT 73.360 199.335 73.500 199.535 ;
        RECT 75.570 199.335 75.890 199.395 ;
        RECT 73.360 199.195 75.890 199.335 ;
        RECT 77.040 199.335 77.180 199.535 ;
        RECT 80.260 199.395 80.400 199.535 ;
        RECT 82.930 199.475 83.250 199.735 ;
        RECT 83.480 199.675 83.620 199.830 ;
        RECT 83.850 199.815 84.170 200.075 ;
        RECT 84.860 200.015 85.000 200.170 ;
        RECT 85.230 200.155 85.550 200.415 ;
        RECT 87.545 200.355 87.835 200.400 ;
        RECT 87.990 200.355 88.310 200.415 ;
        RECT 87.545 200.215 88.310 200.355 ;
        RECT 87.545 200.170 87.835 200.215 ;
        RECT 87.990 200.155 88.310 200.215 ;
        RECT 88.910 200.400 89.230 200.415 ;
        RECT 89.920 200.400 90.060 200.555 ;
        RECT 90.290 200.495 90.610 200.555 ;
        RECT 93.065 200.510 93.355 200.555 ;
        RECT 95.810 200.495 96.130 200.555 ;
        RECT 98.585 200.510 98.875 200.740 ;
        RECT 100.410 200.695 100.730 200.755 ;
        RECT 102.250 200.695 102.570 200.755 ;
        RECT 103.630 200.695 103.950 200.755 ;
        RECT 100.410 200.555 102.570 200.695 ;
        RECT 100.410 200.495 100.730 200.555 ;
        RECT 102.250 200.495 102.570 200.555 ;
        RECT 102.800 200.555 103.950 200.695 ;
        RECT 88.910 200.170 89.365 200.400 ;
        RECT 89.845 200.170 90.135 200.400 ;
        RECT 88.910 200.155 89.230 200.170 ;
        RECT 92.590 200.155 92.910 200.415 ;
        RECT 93.525 200.170 93.815 200.400 ;
        RECT 93.985 200.355 94.275 200.400 ;
        RECT 94.890 200.355 95.210 200.415 ;
        RECT 93.985 200.215 95.210 200.355 ;
        RECT 93.985 200.170 94.275 200.215 ;
        RECT 91.685 200.015 91.975 200.060 ;
        RECT 84.860 199.875 91.975 200.015 ;
        RECT 91.685 199.830 91.975 199.875 ;
        RECT 93.050 200.015 93.370 200.075 ;
        RECT 93.600 200.015 93.740 200.170 ;
        RECT 94.890 200.155 95.210 200.215 ;
        RECT 96.730 200.355 97.050 200.415 ;
        RECT 97.205 200.355 97.495 200.400 ;
        RECT 96.730 200.215 97.495 200.355 ;
        RECT 96.730 200.155 97.050 200.215 ;
        RECT 97.205 200.170 97.495 200.215 ;
        RECT 98.125 200.170 98.415 200.400 ;
        RECT 99.030 200.355 99.350 200.415 ;
        RECT 99.030 200.215 101.100 200.355 ;
        RECT 93.050 199.875 93.740 200.015 ;
        RECT 98.200 200.015 98.340 200.170 ;
        RECT 99.030 200.155 99.350 200.215 ;
        RECT 100.410 200.015 100.730 200.075 ;
        RECT 98.200 199.875 100.730 200.015 ;
        RECT 93.050 199.815 93.370 199.875 ;
        RECT 86.625 199.675 86.915 199.720 ;
        RECT 88.005 199.675 88.295 199.720 ;
        RECT 83.480 199.535 88.295 199.675 ;
        RECT 86.625 199.490 86.915 199.535 ;
        RECT 88.005 199.490 88.295 199.535 ;
        RECT 96.730 199.675 97.050 199.735 ;
        RECT 98.200 199.675 98.340 199.875 ;
        RECT 100.410 199.815 100.730 199.875 ;
        RECT 96.730 199.535 98.340 199.675 ;
        RECT 100.960 199.675 101.100 200.215 ;
        RECT 101.790 200.155 102.110 200.415 ;
        RECT 102.800 200.400 102.940 200.555 ;
        RECT 103.630 200.495 103.950 200.555 ;
        RECT 105.945 200.695 106.235 200.740 ;
        RECT 107.400 200.695 107.540 200.895 ;
        RECT 109.150 200.835 109.470 200.895 ;
        RECT 120.280 200.895 122.350 201.035 ;
        RECT 105.945 200.555 107.540 200.695 ;
        RECT 105.945 200.510 106.235 200.555 ;
        RECT 107.770 200.495 108.090 200.755 ;
        RECT 116.065 200.695 116.355 200.740 ;
        RECT 120.280 200.695 120.420 200.895 ;
        RECT 122.030 200.835 122.350 200.895 ;
        RECT 124.790 200.835 125.110 201.095 ;
        RECT 126.185 201.035 126.475 201.080 ;
        RECT 130.770 201.035 131.090 201.095 ;
        RECT 126.185 200.895 131.090 201.035 ;
        RECT 126.185 200.850 126.475 200.895 ;
        RECT 130.770 200.835 131.090 200.895 ;
        RECT 133.070 201.035 133.390 201.095 ;
        RECT 141.350 201.035 141.670 201.095 ;
        RECT 133.070 200.895 141.670 201.035 ;
        RECT 133.070 200.835 133.390 200.895 ;
        RECT 141.350 200.835 141.670 200.895 ;
        RECT 116.065 200.555 120.420 200.695 ;
        RECT 121.110 200.695 121.430 200.755 ;
        RECT 129.390 200.695 129.710 200.755 ;
        RECT 121.110 200.555 124.100 200.695 ;
        RECT 116.065 200.510 116.355 200.555 ;
        RECT 121.110 200.495 121.430 200.555 ;
        RECT 102.725 200.170 103.015 200.400 ;
        RECT 103.170 200.155 103.490 200.415 ;
        RECT 104.090 200.400 104.410 200.415 ;
        RECT 104.070 200.355 104.410 200.400 ;
        RECT 103.895 200.215 104.410 200.355 ;
        RECT 104.070 200.170 104.410 200.215 ;
        RECT 104.090 200.155 104.410 200.170 ;
        RECT 104.550 200.400 104.870 200.415 ;
        RECT 104.550 200.170 105.085 200.400 ;
        RECT 104.550 200.155 104.870 200.170 ;
        RECT 105.470 200.155 105.790 200.415 ;
        RECT 106.405 200.355 106.695 200.400 ;
        RECT 116.510 200.355 116.830 200.415 ;
        RECT 106.020 200.215 116.830 200.355 ;
        RECT 101.330 200.015 101.650 200.075 ;
        RECT 102.265 200.015 102.555 200.060 ;
        RECT 106.020 200.015 106.160 200.215 ;
        RECT 106.405 200.170 106.695 200.215 ;
        RECT 116.510 200.155 116.830 200.215 ;
        RECT 118.350 200.155 118.670 200.415 ;
        RECT 121.585 200.355 121.875 200.400 ;
        RECT 122.045 200.355 122.335 200.400 ;
        RECT 121.585 200.215 122.335 200.355 ;
        RECT 121.585 200.170 121.875 200.215 ;
        RECT 122.045 200.170 122.335 200.215 ;
        RECT 122.965 200.170 123.255 200.400 ;
        RECT 115.590 200.015 115.910 200.075 ;
        RECT 101.330 199.875 102.555 200.015 ;
        RECT 101.330 199.815 101.650 199.875 ;
        RECT 102.265 199.830 102.555 199.875 ;
        RECT 104.640 199.875 106.160 200.015 ;
        RECT 106.480 199.875 115.910 200.015 ;
        RECT 104.640 199.675 104.780 199.875 ;
        RECT 100.960 199.535 104.780 199.675 ;
        RECT 105.010 199.675 105.330 199.735 ;
        RECT 106.480 199.675 106.620 199.875 ;
        RECT 115.590 199.815 115.910 199.875 ;
        RECT 116.050 200.015 116.370 200.075 ;
        RECT 121.110 200.015 121.430 200.075 ;
        RECT 116.050 199.875 121.430 200.015 ;
        RECT 123.040 200.015 123.180 200.170 ;
        RECT 123.410 200.155 123.730 200.415 ;
        RECT 123.960 200.400 124.100 200.555 ;
        RECT 126.720 200.555 129.710 200.695 ;
        RECT 123.885 200.170 124.175 200.400 ;
        RECT 126.720 200.015 126.860 200.555 ;
        RECT 129.390 200.495 129.710 200.555 ;
        RECT 129.850 200.695 130.170 200.755 ;
        RECT 129.850 200.555 139.740 200.695 ;
        RECT 129.850 200.495 130.170 200.555 ;
        RECT 127.550 200.155 127.870 200.415 ;
        RECT 128.930 200.155 129.250 200.415 ;
        RECT 134.910 200.355 135.230 200.415 ;
        RECT 136.290 200.355 136.610 200.415 ;
        RECT 129.480 200.215 136.610 200.355 ;
        RECT 129.480 200.060 129.620 200.215 ;
        RECT 134.910 200.155 135.230 200.215 ;
        RECT 136.290 200.155 136.610 200.215 ;
        RECT 137.210 200.155 137.530 200.415 ;
        RECT 138.605 200.355 138.895 200.400 ;
        RECT 139.050 200.355 139.370 200.415 ;
        RECT 139.600 200.400 139.740 200.555 ;
        RECT 138.605 200.215 139.370 200.355 ;
        RECT 138.605 200.170 138.895 200.215 ;
        RECT 139.050 200.155 139.370 200.215 ;
        RECT 139.525 200.170 139.815 200.400 ;
        RECT 140.890 200.155 141.210 200.415 ;
        RECT 143.190 200.155 143.510 200.415 ;
        RECT 144.585 200.170 144.875 200.400 ;
        RECT 123.040 199.875 126.860 200.015 ;
        RECT 116.050 199.815 116.370 199.875 ;
        RECT 121.110 199.815 121.430 199.875 ;
        RECT 127.105 199.830 127.395 200.060 ;
        RECT 129.405 199.830 129.695 200.060 ;
        RECT 105.010 199.535 106.620 199.675 ;
        RECT 110.530 199.675 110.850 199.735 ;
        RECT 126.170 199.675 126.490 199.735 ;
        RECT 127.180 199.675 127.320 199.830 ;
        RECT 133.530 199.815 133.850 200.075 ;
        RECT 134.450 199.815 134.770 200.075 ;
        RECT 144.660 200.015 144.800 200.170 ;
        RECT 135.460 199.875 144.800 200.015 ;
        RECT 135.460 199.675 135.600 199.875 ;
        RECT 110.530 199.535 125.940 199.675 ;
        RECT 96.730 199.475 97.050 199.535 ;
        RECT 105.010 199.475 105.330 199.535 ;
        RECT 110.530 199.475 110.850 199.535 ;
        RECT 78.790 199.335 79.110 199.395 ;
        RECT 77.040 199.195 79.110 199.335 ;
        RECT 36.470 199.135 36.790 199.195 ;
        RECT 41.530 199.135 41.850 199.195 ;
        RECT 47.970 199.135 48.290 199.195 ;
        RECT 51.205 199.150 51.495 199.195 ;
        RECT 56.250 199.135 56.570 199.195 ;
        RECT 71.445 199.150 71.735 199.195 ;
        RECT 75.570 199.135 75.890 199.195 ;
        RECT 78.790 199.135 79.110 199.195 ;
        RECT 80.170 199.135 80.490 199.395 ;
        RECT 86.150 199.380 86.470 199.395 ;
        RECT 85.935 199.150 86.470 199.380 ;
        RECT 86.150 199.135 86.470 199.150 ;
        RECT 87.070 199.135 87.390 199.395 ;
        RECT 94.430 199.335 94.750 199.395 ;
        RECT 99.030 199.335 99.350 199.395 ;
        RECT 94.430 199.195 99.350 199.335 ;
        RECT 94.430 199.135 94.750 199.195 ;
        RECT 99.030 199.135 99.350 199.195 ;
        RECT 99.965 199.335 100.255 199.380 ;
        RECT 100.870 199.335 101.190 199.395 ;
        RECT 99.965 199.195 101.190 199.335 ;
        RECT 99.965 199.150 100.255 199.195 ;
        RECT 100.870 199.135 101.190 199.195 ;
        RECT 102.710 199.335 103.030 199.395 ;
        RECT 103.645 199.335 103.935 199.380 ;
        RECT 102.710 199.195 103.935 199.335 ;
        RECT 102.710 199.135 103.030 199.195 ;
        RECT 103.645 199.150 103.935 199.195 ;
        RECT 107.310 199.135 107.630 199.395 ;
        RECT 111.450 199.335 111.770 199.395 ;
        RECT 123.410 199.335 123.730 199.395 ;
        RECT 111.450 199.195 123.730 199.335 ;
        RECT 125.800 199.335 125.940 199.535 ;
        RECT 126.170 199.535 127.320 199.675 ;
        RECT 127.640 199.535 135.600 199.675 ;
        RECT 135.845 199.675 136.135 199.720 ;
        RECT 138.605 199.675 138.895 199.720 ;
        RECT 139.510 199.675 139.830 199.735 ;
        RECT 135.845 199.535 138.360 199.675 ;
        RECT 126.170 199.475 126.490 199.535 ;
        RECT 127.640 199.335 127.780 199.535 ;
        RECT 135.845 199.490 136.135 199.535 ;
        RECT 125.800 199.195 127.780 199.335 ;
        RECT 128.010 199.335 128.330 199.395 ;
        RECT 130.785 199.335 131.075 199.380 ;
        RECT 128.010 199.195 131.075 199.335 ;
        RECT 111.450 199.135 111.770 199.195 ;
        RECT 123.410 199.135 123.730 199.195 ;
        RECT 128.010 199.135 128.330 199.195 ;
        RECT 130.785 199.150 131.075 199.195 ;
        RECT 131.690 199.335 132.010 199.395 ;
        RECT 135.920 199.335 136.060 199.490 ;
        RECT 131.690 199.195 136.060 199.335 ;
        RECT 131.690 199.135 132.010 199.195 ;
        RECT 136.750 199.135 137.070 199.395 ;
        RECT 137.210 199.335 137.530 199.395 ;
        RECT 137.685 199.335 137.975 199.380 ;
        RECT 137.210 199.195 137.975 199.335 ;
        RECT 138.220 199.335 138.360 199.535 ;
        RECT 138.605 199.535 139.830 199.675 ;
        RECT 138.605 199.490 138.895 199.535 ;
        RECT 139.510 199.475 139.830 199.535 ;
        RECT 145.490 199.475 145.810 199.735 ;
        RECT 139.050 199.335 139.370 199.395 ;
        RECT 138.220 199.195 139.370 199.335 ;
        RECT 137.210 199.135 137.530 199.195 ;
        RECT 137.685 199.150 137.975 199.195 ;
        RECT 139.050 199.135 139.370 199.195 ;
        RECT 141.810 199.135 142.130 199.395 ;
        RECT 143.650 199.135 143.970 199.395 ;
        RECT 13.860 198.515 147.720 198.995 ;
        RECT 14.850 198.315 15.170 198.375 ;
        RECT 15.785 198.315 16.075 198.360 ;
        RECT 14.850 198.175 16.075 198.315 ;
        RECT 14.850 198.115 15.170 198.175 ;
        RECT 15.785 198.130 16.075 198.175 ;
        RECT 28.190 198.315 28.510 198.375 ;
        RECT 30.490 198.315 30.810 198.375 ;
        RECT 28.190 198.175 30.810 198.315 ;
        RECT 28.190 198.115 28.510 198.175 ;
        RECT 30.490 198.115 30.810 198.175 ;
        RECT 35.090 198.315 35.410 198.375 ;
        RECT 36.470 198.315 36.790 198.375 ;
        RECT 35.090 198.175 36.790 198.315 ;
        RECT 35.090 198.115 35.410 198.175 ;
        RECT 36.470 198.115 36.790 198.175 ;
        RECT 36.930 198.315 37.250 198.375 ;
        RECT 38.325 198.315 38.615 198.360 ;
        RECT 36.930 198.175 38.615 198.315 ;
        RECT 36.930 198.115 37.250 198.175 ;
        RECT 38.325 198.130 38.615 198.175 ;
        RECT 39.230 198.115 39.550 198.375 ;
        RECT 40.610 198.315 40.930 198.375 ;
        RECT 42.005 198.315 42.295 198.360 ;
        RECT 40.610 198.175 42.295 198.315 ;
        RECT 40.610 198.115 40.930 198.175 ;
        RECT 42.005 198.130 42.295 198.175 ;
        RECT 48.890 198.315 49.210 198.375 ;
        RECT 51.650 198.315 51.970 198.375 ;
        RECT 48.890 198.175 51.970 198.315 ;
        RECT 48.890 198.115 49.210 198.175 ;
        RECT 51.650 198.115 51.970 198.175 ;
        RECT 54.870 198.315 55.190 198.375 ;
        RECT 58.090 198.315 58.410 198.375 ;
        RECT 54.870 198.175 58.410 198.315 ;
        RECT 54.870 198.115 55.190 198.175 ;
        RECT 58.090 198.115 58.410 198.175 ;
        RECT 58.550 198.315 58.870 198.375 ;
        RECT 59.025 198.315 59.315 198.360 ;
        RECT 58.550 198.175 59.315 198.315 ;
        RECT 58.550 198.115 58.870 198.175 ;
        RECT 59.025 198.130 59.315 198.175 ;
        RECT 63.150 198.315 63.470 198.375 ;
        RECT 71.430 198.315 71.750 198.375 ;
        RECT 74.665 198.315 74.955 198.360 ;
        RECT 63.150 198.175 74.955 198.315 ;
        RECT 63.150 198.115 63.470 198.175 ;
        RECT 71.430 198.115 71.750 198.175 ;
        RECT 74.665 198.130 74.955 198.175 ;
        RECT 82.945 198.315 83.235 198.360 ;
        RECT 83.390 198.315 83.710 198.375 ;
        RECT 82.945 198.175 83.710 198.315 ;
        RECT 82.945 198.130 83.235 198.175 ;
        RECT 83.390 198.115 83.710 198.175 ;
        RECT 97.650 198.115 97.970 198.375 ;
        RECT 103.645 198.315 103.935 198.360 ;
        RECT 105.470 198.315 105.790 198.375 ;
        RECT 103.645 198.175 105.790 198.315 ;
        RECT 103.645 198.130 103.935 198.175 ;
        RECT 105.470 198.115 105.790 198.175 ;
        RECT 109.610 198.115 109.930 198.375 ;
        RECT 127.550 198.315 127.870 198.375 ;
        RECT 139.510 198.315 139.830 198.375 ;
        RECT 111.540 198.175 127.870 198.315 ;
        RECT 18.495 197.975 18.785 198.020 ;
        RECT 20.385 197.975 20.675 198.020 ;
        RECT 23.505 197.975 23.795 198.020 ;
        RECT 18.495 197.835 23.795 197.975 ;
        RECT 18.495 197.790 18.785 197.835 ;
        RECT 20.385 197.790 20.675 197.835 ;
        RECT 23.505 197.790 23.795 197.835 ;
        RECT 24.510 197.975 24.830 198.035 ;
        RECT 25.890 197.975 26.210 198.035 ;
        RECT 24.510 197.835 26.210 197.975 ;
        RECT 24.510 197.775 24.830 197.835 ;
        RECT 25.890 197.775 26.210 197.835 ;
        RECT 32.790 197.975 33.110 198.035 ;
        RECT 34.630 197.975 34.950 198.035 ;
        RECT 60.815 197.975 61.105 198.020 ;
        RECT 62.705 197.975 62.995 198.020 ;
        RECT 65.825 197.975 66.115 198.020 ;
        RECT 32.790 197.835 33.940 197.975 ;
        RECT 32.790 197.775 33.110 197.835 ;
        RECT 17.625 197.635 17.915 197.680 ;
        RECT 18.990 197.635 19.310 197.695 ;
        RECT 17.625 197.495 19.310 197.635 ;
        RECT 17.625 197.450 17.915 197.495 ;
        RECT 18.990 197.435 19.310 197.495 ;
        RECT 22.210 197.635 22.530 197.695 ;
        RECT 26.365 197.635 26.655 197.680 ;
        RECT 32.330 197.635 32.650 197.695 ;
        RECT 22.210 197.495 26.120 197.635 ;
        RECT 22.210 197.435 22.530 197.495 ;
        RECT 16.705 197.295 16.995 197.340 ;
        RECT 17.150 197.295 17.470 197.355 ;
        RECT 16.705 197.155 17.470 197.295 ;
        RECT 16.705 197.110 16.995 197.155 ;
        RECT 17.150 197.095 17.470 197.155 ;
        RECT 18.090 197.295 18.380 197.340 ;
        RECT 19.925 197.295 20.215 197.340 ;
        RECT 23.505 197.295 23.795 197.340 ;
        RECT 18.090 197.155 23.795 197.295 ;
        RECT 18.090 197.110 18.380 197.155 ;
        RECT 19.925 197.110 20.215 197.155 ;
        RECT 23.505 197.110 23.795 197.155 ;
        RECT 24.510 197.315 24.830 197.355 ;
        RECT 24.510 197.095 24.875 197.315 ;
        RECT 25.980 197.295 26.120 197.495 ;
        RECT 26.365 197.495 32.650 197.635 ;
        RECT 26.365 197.450 26.655 197.495 ;
        RECT 28.205 197.295 28.495 197.340 ;
        RECT 28.650 197.295 28.970 197.355 ;
        RECT 25.980 197.155 28.970 197.295 ;
        RECT 28.205 197.110 28.495 197.155 ;
        RECT 28.650 197.095 28.970 197.155 ;
        RECT 29.585 197.295 29.875 197.340 ;
        RECT 30.030 197.295 30.350 197.355 ;
        RECT 31.500 197.340 31.640 197.495 ;
        RECT 32.330 197.435 32.650 197.495 ;
        RECT 29.585 197.155 30.350 197.295 ;
        RECT 29.585 197.110 29.875 197.155 ;
        RECT 30.030 197.095 30.350 197.155 ;
        RECT 31.425 197.110 31.715 197.340 ;
        RECT 31.885 197.110 32.175 197.340 ;
        RECT 32.805 197.110 33.095 197.340 ;
        RECT 24.585 197.000 24.875 197.095 ;
        RECT 19.005 196.770 19.295 197.000 ;
        RECT 21.285 196.955 21.935 197.000 ;
        RECT 24.585 196.955 25.175 197.000 ;
        RECT 27.285 196.955 27.575 197.000 ;
        RECT 31.960 196.955 32.100 197.110 ;
        RECT 21.285 196.815 25.175 196.955 ;
        RECT 21.285 196.770 21.935 196.815 ;
        RECT 24.885 196.770 25.175 196.815 ;
        RECT 25.520 196.815 27.575 196.955 ;
        RECT 19.080 196.615 19.220 196.770 ;
        RECT 25.520 196.615 25.660 196.815 ;
        RECT 27.285 196.770 27.575 196.815 ;
        RECT 31.500 196.815 32.100 196.955 ;
        RECT 32.880 196.955 33.020 197.110 ;
        RECT 33.250 197.095 33.570 197.355 ;
        RECT 33.800 197.340 33.940 197.835 ;
        RECT 34.630 197.835 57.860 197.975 ;
        RECT 34.630 197.775 34.950 197.835 ;
        RECT 35.105 197.635 35.395 197.680 ;
        RECT 38.310 197.635 38.630 197.695 ;
        RECT 35.105 197.495 36.700 197.635 ;
        RECT 35.105 197.450 35.395 197.495 ;
        RECT 33.725 197.295 34.015 197.340 ;
        RECT 35.550 197.295 35.870 197.355 ;
        RECT 36.560 197.340 36.700 197.495 ;
        RECT 37.480 197.495 38.630 197.635 ;
        RECT 33.725 197.155 35.870 197.295 ;
        RECT 33.725 197.110 34.015 197.155 ;
        RECT 35.550 197.095 35.870 197.155 ;
        RECT 36.485 197.110 36.775 197.340 ;
        RECT 37.480 196.955 37.620 197.495 ;
        RECT 38.310 197.435 38.630 197.495 ;
        RECT 39.705 197.635 39.995 197.680 ;
        RECT 41.070 197.635 41.390 197.695 ;
        RECT 39.705 197.495 41.390 197.635 ;
        RECT 39.705 197.450 39.995 197.495 ;
        RECT 41.070 197.435 41.390 197.495 ;
        RECT 43.370 197.635 43.690 197.695 ;
        RECT 43.370 197.495 44.980 197.635 ;
        RECT 43.370 197.435 43.690 197.495 ;
        RECT 37.865 197.110 38.155 197.340 ;
        RECT 32.880 196.815 37.620 196.955 ;
        RECT 37.940 196.955 38.080 197.110 ;
        RECT 40.150 197.095 40.470 197.355 ;
        RECT 41.545 197.110 41.835 197.340 ;
        RECT 42.465 197.295 42.755 197.340 ;
        RECT 42.910 197.295 43.230 197.355 ;
        RECT 44.840 197.340 44.980 197.495 ;
        RECT 48.890 197.435 49.210 197.695 ;
        RECT 50.730 197.635 51.050 197.695 ;
        RECT 56.250 197.635 56.570 197.695 ;
        RECT 57.720 197.635 57.860 197.835 ;
        RECT 60.815 197.835 66.115 197.975 ;
        RECT 60.815 197.790 61.105 197.835 ;
        RECT 62.705 197.790 62.995 197.835 ;
        RECT 65.825 197.790 66.115 197.835 ;
        RECT 66.830 197.975 67.150 198.035 ;
        RECT 68.210 197.975 68.530 198.035 ;
        RECT 72.350 197.975 72.670 198.035 ;
        RECT 66.830 197.835 68.530 197.975 ;
        RECT 66.830 197.775 67.150 197.835 ;
        RECT 68.210 197.775 68.530 197.835 ;
        RECT 69.220 197.835 72.670 197.975 ;
        RECT 59.945 197.635 60.235 197.680 ;
        RECT 66.920 197.635 67.060 197.775 ;
        RECT 50.730 197.495 54.180 197.635 ;
        RECT 50.730 197.435 51.050 197.495 ;
        RECT 43.845 197.295 44.135 197.340 ;
        RECT 42.465 197.155 44.135 197.295 ;
        RECT 42.465 197.110 42.755 197.155 ;
        RECT 39.230 196.955 39.550 197.015 ;
        RECT 41.620 196.955 41.760 197.110 ;
        RECT 42.910 197.095 43.230 197.155 ;
        RECT 43.845 197.110 44.135 197.155 ;
        RECT 44.765 197.110 45.055 197.340 ;
        RECT 45.670 197.295 45.990 197.355 ;
        RECT 47.985 197.295 48.275 197.340 ;
        RECT 49.825 197.295 50.115 197.340 ;
        RECT 45.670 197.155 48.275 197.295 ;
        RECT 45.670 197.095 45.990 197.155 ;
        RECT 47.985 197.110 48.275 197.155 ;
        RECT 48.980 197.155 50.115 197.295 ;
        RECT 37.940 196.815 41.760 196.955 ;
        RECT 31.500 196.675 31.640 196.815 ;
        RECT 39.230 196.755 39.550 196.815 ;
        RECT 46.145 196.770 46.435 197.000 ;
        RECT 46.605 196.955 46.895 197.000 ;
        RECT 47.050 196.955 47.370 197.015 ;
        RECT 48.980 196.955 49.120 197.155 ;
        RECT 49.825 197.110 50.115 197.155 ;
        RECT 50.285 197.110 50.575 197.340 ;
        RECT 51.205 197.295 51.495 197.340 ;
        RECT 51.650 197.295 51.970 197.355 ;
        RECT 53.030 197.295 53.350 197.355 ;
        RECT 54.040 197.340 54.180 197.495 ;
        RECT 56.250 197.495 57.400 197.635 ;
        RECT 57.720 197.495 59.240 197.635 ;
        RECT 56.250 197.435 56.570 197.495 ;
        RECT 57.260 197.340 57.400 197.495 ;
        RECT 59.100 197.355 59.240 197.495 ;
        RECT 59.945 197.495 67.060 197.635 ;
        RECT 59.945 197.450 60.235 197.495 ;
        RECT 51.205 197.155 51.970 197.295 ;
        RECT 51.205 197.110 51.495 197.155 ;
        RECT 46.605 196.815 49.120 196.955 ;
        RECT 46.605 196.770 46.895 196.815 ;
        RECT 19.080 196.475 25.660 196.615 ;
        RECT 26.350 196.615 26.670 196.675 ;
        RECT 28.190 196.615 28.510 196.675 ;
        RECT 29.125 196.615 29.415 196.660 ;
        RECT 30.505 196.615 30.795 196.660 ;
        RECT 26.350 196.475 30.795 196.615 ;
        RECT 26.350 196.415 26.670 196.475 ;
        RECT 28.190 196.415 28.510 196.475 ;
        RECT 29.125 196.430 29.415 196.475 ;
        RECT 30.505 196.430 30.795 196.475 ;
        RECT 31.410 196.415 31.730 196.675 ;
        RECT 32.330 196.615 32.650 196.675 ;
        RECT 35.565 196.615 35.855 196.660 ;
        RECT 32.330 196.475 35.855 196.615 ;
        RECT 32.330 196.415 32.650 196.475 ;
        RECT 35.565 196.430 35.855 196.475 ;
        RECT 37.405 196.615 37.695 196.660 ;
        RECT 42.910 196.615 43.230 196.675 ;
        RECT 37.405 196.475 43.230 196.615 ;
        RECT 46.220 196.615 46.360 196.770 ;
        RECT 47.050 196.755 47.370 196.815 ;
        RECT 49.350 196.755 49.670 197.015 ;
        RECT 50.360 196.955 50.500 197.110 ;
        RECT 51.650 197.095 51.970 197.155 ;
        RECT 52.660 197.155 53.350 197.295 ;
        RECT 52.110 196.955 52.430 197.015 ;
        RECT 50.360 196.815 52.430 196.955 ;
        RECT 52.110 196.755 52.430 196.815 ;
        RECT 48.890 196.615 49.210 196.675 ;
        RECT 46.220 196.475 49.210 196.615 ;
        RECT 37.405 196.430 37.695 196.475 ;
        RECT 42.910 196.415 43.230 196.475 ;
        RECT 48.890 196.415 49.210 196.475 ;
        RECT 50.745 196.615 51.035 196.660 ;
        RECT 52.660 196.615 52.800 197.155 ;
        RECT 53.030 197.095 53.350 197.155 ;
        RECT 53.965 197.110 54.255 197.340 ;
        RECT 56.725 197.110 57.015 197.340 ;
        RECT 57.185 197.110 57.475 197.340 ;
        RECT 56.800 196.955 56.940 197.110 ;
        RECT 58.090 197.095 58.410 197.355 ;
        RECT 58.565 197.110 58.855 197.340 ;
        RECT 58.180 196.955 58.320 197.095 ;
        RECT 56.800 196.815 58.320 196.955 ;
        RECT 50.745 196.475 52.800 196.615 ;
        RECT 50.745 196.430 51.035 196.475 ;
        RECT 53.030 196.415 53.350 196.675 ;
        RECT 55.330 196.615 55.650 196.675 ;
        RECT 56.265 196.615 56.555 196.660 ;
        RECT 55.330 196.475 56.555 196.615 ;
        RECT 55.330 196.415 55.650 196.475 ;
        RECT 56.265 196.430 56.555 196.475 ;
        RECT 57.630 196.415 57.950 196.675 ;
        RECT 58.090 196.615 58.410 196.675 ;
        RECT 58.640 196.615 58.780 197.110 ;
        RECT 59.010 197.095 59.330 197.355 ;
        RECT 59.470 197.095 59.790 197.355 ;
        RECT 60.410 197.295 60.700 197.340 ;
        RECT 62.245 197.295 62.535 197.340 ;
        RECT 65.825 197.295 66.115 197.340 ;
        RECT 60.410 197.155 66.115 197.295 ;
        RECT 60.410 197.110 60.700 197.155 ;
        RECT 62.245 197.110 62.535 197.155 ;
        RECT 65.825 197.110 66.115 197.155 ;
        RECT 66.370 197.295 66.690 197.355 ;
        RECT 66.905 197.295 67.195 197.315 ;
        RECT 68.670 197.295 68.990 197.355 ;
        RECT 66.370 197.155 68.990 197.295 ;
        RECT 66.370 197.095 66.690 197.155 ;
        RECT 61.310 196.755 61.630 197.015 ;
        RECT 66.905 197.000 67.195 197.155 ;
        RECT 68.670 197.095 68.990 197.155 ;
        RECT 63.605 196.955 64.255 197.000 ;
        RECT 66.905 196.955 67.495 197.000 ;
        RECT 69.220 196.955 69.360 197.835 ;
        RECT 72.350 197.775 72.670 197.835 ;
        RECT 75.585 197.975 75.875 198.020 ;
        RECT 97.190 197.975 97.510 198.035 ;
        RECT 75.585 197.835 97.510 197.975 ;
        RECT 75.585 197.790 75.875 197.835 ;
        RECT 97.190 197.775 97.510 197.835 ;
        RECT 70.065 197.635 70.355 197.680 ;
        RECT 71.430 197.635 71.750 197.695 ;
        RECT 73.270 197.635 73.590 197.695 ;
        RECT 74.190 197.635 74.510 197.695 ;
        RECT 70.065 197.495 71.750 197.635 ;
        RECT 70.065 197.450 70.355 197.495 ;
        RECT 71.430 197.435 71.750 197.495 ;
        RECT 71.980 197.495 74.510 197.635 ;
        RECT 69.590 197.295 69.910 197.355 ;
        RECT 70.525 197.295 70.815 197.340 ;
        RECT 71.980 197.295 72.120 197.495 ;
        RECT 73.270 197.435 73.590 197.495 ;
        RECT 74.190 197.435 74.510 197.495 ;
        RECT 74.650 197.635 74.970 197.695 ;
        RECT 83.865 197.635 84.155 197.680 ;
        RECT 86.150 197.635 86.470 197.695 ;
        RECT 95.350 197.635 95.670 197.695 ;
        RECT 74.650 197.495 81.320 197.635 ;
        RECT 74.650 197.435 74.970 197.495 ;
        RECT 69.590 197.155 72.120 197.295 ;
        RECT 72.350 197.295 72.670 197.355 ;
        RECT 72.350 197.155 77.180 197.295 ;
        RECT 69.590 197.095 69.910 197.155 ;
        RECT 70.525 197.110 70.815 197.155 ;
        RECT 72.350 197.095 72.670 197.155 ;
        RECT 63.605 196.815 67.495 196.955 ;
        RECT 63.605 196.770 64.255 196.815 ;
        RECT 67.205 196.770 67.495 196.815 ;
        RECT 67.840 196.815 69.360 196.955 ;
        RECT 67.840 196.615 67.980 196.815 ;
        RECT 58.090 196.475 67.980 196.615 ;
        RECT 68.210 196.615 68.530 196.675 ;
        RECT 69.680 196.615 69.820 197.095 ;
        RECT 73.730 196.955 74.050 197.015 ;
        RECT 73.730 196.815 75.340 196.955 ;
        RECT 73.730 196.755 74.050 196.815 ;
        RECT 68.210 196.475 69.820 196.615 ;
        RECT 58.090 196.415 58.410 196.475 ;
        RECT 68.210 196.415 68.530 196.475 ;
        RECT 71.430 196.415 71.750 196.675 ;
        RECT 71.890 196.415 72.210 196.675 ;
        RECT 72.365 196.615 72.655 196.660 ;
        RECT 72.810 196.615 73.130 196.675 ;
        RECT 72.365 196.475 73.130 196.615 ;
        RECT 72.365 196.430 72.655 196.475 ;
        RECT 72.810 196.415 73.130 196.475 ;
        RECT 73.270 196.415 73.590 196.675 ;
        RECT 74.650 196.660 74.970 196.675 ;
        RECT 74.650 196.430 75.035 196.660 ;
        RECT 75.200 196.615 75.340 196.815 ;
        RECT 76.490 196.615 76.810 196.675 ;
        RECT 77.040 196.660 77.180 197.155 ;
        RECT 77.870 197.095 78.190 197.355 ;
        RECT 78.790 197.095 79.110 197.355 ;
        RECT 80.630 197.095 80.950 197.355 ;
        RECT 79.710 196.755 80.030 197.015 ;
        RECT 80.185 196.770 80.475 197.000 ;
        RECT 81.180 196.955 81.320 197.495 ;
        RECT 83.865 197.495 86.470 197.635 ;
        RECT 83.865 197.450 84.155 197.495 ;
        RECT 86.150 197.435 86.470 197.495 ;
        RECT 86.700 197.495 95.670 197.635 ;
        RECT 97.740 197.635 97.880 198.115 ;
        RECT 98.570 197.975 98.890 198.035 ;
        RECT 104.090 197.975 104.410 198.035 ;
        RECT 98.570 197.835 104.410 197.975 ;
        RECT 98.570 197.775 98.890 197.835 ;
        RECT 104.090 197.775 104.410 197.835 ;
        RECT 104.550 197.975 104.870 198.035 ;
        RECT 106.390 197.975 106.710 198.035 ;
        RECT 104.550 197.835 106.710 197.975 ;
        RECT 104.550 197.775 104.870 197.835 ;
        RECT 106.390 197.775 106.710 197.835 ;
        RECT 107.325 197.975 107.615 198.020 ;
        RECT 111.540 197.975 111.680 198.175 ;
        RECT 127.550 198.115 127.870 198.175 ;
        RECT 132.240 198.175 139.830 198.315 ;
        RECT 107.325 197.835 111.680 197.975 ;
        RECT 111.875 197.975 112.165 198.020 ;
        RECT 113.765 197.975 114.055 198.020 ;
        RECT 116.885 197.975 117.175 198.020 ;
        RECT 111.875 197.835 117.175 197.975 ;
        RECT 107.325 197.790 107.615 197.835 ;
        RECT 111.875 197.790 112.165 197.835 ;
        RECT 113.765 197.790 114.055 197.835 ;
        RECT 116.885 197.790 117.175 197.835 ;
        RECT 123.410 197.975 123.730 198.035 ;
        RECT 125.725 197.975 126.015 198.020 ;
        RECT 123.410 197.835 131.460 197.975 ;
        RECT 123.410 197.775 123.730 197.835 ;
        RECT 125.725 197.790 126.015 197.835 ;
        RECT 98.125 197.635 98.415 197.680 ;
        RECT 97.740 197.495 98.415 197.635 ;
        RECT 84.310 197.095 84.630 197.355 ;
        RECT 84.770 197.095 85.090 197.355 ;
        RECT 86.700 196.955 86.840 197.495 ;
        RECT 95.350 197.435 95.670 197.495 ;
        RECT 98.125 197.450 98.415 197.495 ;
        RECT 100.410 197.635 100.730 197.695 ;
        RECT 107.785 197.635 108.075 197.680 ;
        RECT 108.690 197.635 109.010 197.695 ;
        RECT 100.410 197.495 106.620 197.635 ;
        RECT 100.410 197.435 100.730 197.495 ;
        RECT 90.765 197.110 91.055 197.340 ;
        RECT 81.180 196.815 86.840 196.955 ;
        RECT 87.990 196.955 88.310 197.015 ;
        RECT 89.830 196.955 90.150 197.015 ;
        RECT 90.840 196.955 90.980 197.110 ;
        RECT 91.670 197.095 91.990 197.355 ;
        RECT 96.270 197.295 96.590 197.355 ;
        RECT 101.805 197.295 102.095 197.340 ;
        RECT 96.270 197.155 99.260 197.295 ;
        RECT 96.270 197.095 96.590 197.155 ;
        RECT 99.120 197.015 99.260 197.155 ;
        RECT 100.500 197.155 102.095 197.295 ;
        RECT 93.050 196.955 93.370 197.015 ;
        RECT 87.990 196.815 93.370 196.955 ;
        RECT 75.200 196.475 76.810 196.615 ;
        RECT 74.650 196.415 74.970 196.430 ;
        RECT 76.490 196.415 76.810 196.475 ;
        RECT 76.965 196.615 77.255 196.660 ;
        RECT 80.260 196.615 80.400 196.770 ;
        RECT 87.990 196.755 88.310 196.815 ;
        RECT 89.830 196.755 90.150 196.815 ;
        RECT 93.050 196.755 93.370 196.815 ;
        RECT 99.030 196.755 99.350 197.015 ;
        RECT 99.490 196.955 99.810 197.015 ;
        RECT 100.500 196.955 100.640 197.155 ;
        RECT 101.805 197.110 102.095 197.155 ;
        RECT 102.250 197.095 102.570 197.355 ;
        RECT 102.710 197.095 103.030 197.355 ;
        RECT 104.090 197.295 104.410 197.355 ;
        RECT 105.945 197.295 106.235 197.340 ;
        RECT 104.090 197.155 106.235 197.295 ;
        RECT 104.090 197.095 104.410 197.155 ;
        RECT 105.945 197.110 106.235 197.155 ;
        RECT 99.490 196.815 100.640 196.955 ;
        RECT 100.885 196.955 101.175 197.000 ;
        RECT 104.565 196.955 104.855 197.000 ;
        RECT 100.885 196.815 104.855 196.955 ;
        RECT 106.480 196.955 106.620 197.495 ;
        RECT 107.785 197.495 109.010 197.635 ;
        RECT 107.785 197.450 108.075 197.495 ;
        RECT 108.690 197.435 109.010 197.495 ;
        RECT 109.610 197.635 109.930 197.695 ;
        RECT 122.490 197.635 122.810 197.695 ;
        RECT 131.320 197.680 131.460 197.835 ;
        RECT 132.240 197.680 132.380 198.175 ;
        RECT 139.510 198.115 139.830 198.175 ;
        RECT 145.490 198.115 145.810 198.375 ;
        RECT 132.610 197.975 132.930 198.035 ;
        RECT 132.610 197.835 144.800 197.975 ;
        RECT 132.610 197.775 132.930 197.835 ;
        RECT 125.265 197.635 125.555 197.680 ;
        RECT 109.610 197.495 122.260 197.635 ;
        RECT 109.610 197.435 109.930 197.495 ;
        RECT 107.310 197.295 107.630 197.355 ;
        RECT 110.530 197.295 110.850 197.355 ;
        RECT 107.310 197.155 110.850 197.295 ;
        RECT 107.310 197.095 107.630 197.155 ;
        RECT 110.530 197.095 110.850 197.155 ;
        RECT 110.990 197.095 111.310 197.355 ;
        RECT 111.470 197.295 111.760 197.340 ;
        RECT 113.305 197.295 113.595 197.340 ;
        RECT 116.885 197.295 117.175 197.340 ;
        RECT 111.470 197.155 117.175 197.295 ;
        RECT 111.470 197.110 111.760 197.155 ;
        RECT 113.305 197.110 113.595 197.155 ;
        RECT 116.885 197.110 117.175 197.155 ;
        RECT 117.965 197.295 118.255 197.315 ;
        RECT 122.120 197.295 122.260 197.495 ;
        RECT 122.490 197.495 125.555 197.635 ;
        RECT 122.490 197.435 122.810 197.495 ;
        RECT 125.265 197.450 125.555 197.495 ;
        RECT 131.245 197.450 131.535 197.680 ;
        RECT 132.165 197.450 132.455 197.680 ;
        RECT 135.385 197.635 135.675 197.680 ;
        RECT 143.650 197.635 143.970 197.695 ;
        RECT 135.385 197.495 143.970 197.635 ;
        RECT 135.385 197.450 135.675 197.495 ;
        RECT 143.650 197.435 143.970 197.495 ;
        RECT 124.345 197.295 124.635 197.340 ;
        RECT 126.170 197.295 126.490 197.355 ;
        RECT 117.965 197.155 121.800 197.295 ;
        RECT 122.120 197.155 126.490 197.295 ;
        RECT 109.625 196.955 109.915 197.000 ;
        RECT 106.480 196.815 109.915 196.955 ;
        RECT 99.490 196.755 99.810 196.815 ;
        RECT 100.885 196.770 101.175 196.815 ;
        RECT 104.565 196.770 104.855 196.815 ;
        RECT 109.625 196.770 109.915 196.815 ;
        RECT 112.370 196.755 112.690 197.015 ;
        RECT 117.965 197.000 118.255 197.155 ;
        RECT 114.665 196.955 115.315 197.000 ;
        RECT 117.965 196.955 118.555 197.000 ;
        RECT 114.665 196.815 118.555 196.955 ;
        RECT 114.665 196.770 115.315 196.815 ;
        RECT 118.265 196.770 118.555 196.815 ;
        RECT 119.730 196.955 120.050 197.015 ;
        RECT 121.125 196.955 121.415 197.000 ;
        RECT 119.730 196.815 121.415 196.955 ;
        RECT 121.660 196.955 121.800 197.155 ;
        RECT 124.345 197.110 124.635 197.155 ;
        RECT 126.170 197.095 126.490 197.155 ;
        RECT 126.645 197.275 126.935 197.340 ;
        RECT 128.010 197.275 128.330 197.355 ;
        RECT 126.645 197.135 128.330 197.275 ;
        RECT 126.645 197.110 126.935 197.135 ;
        RECT 128.010 197.095 128.330 197.135 ;
        RECT 129.390 197.095 129.710 197.355 ;
        RECT 131.690 197.295 132.010 197.355 ;
        RECT 133.545 197.295 133.835 197.340 ;
        RECT 136.765 197.295 137.055 197.340 ;
        RECT 131.690 197.155 133.835 197.295 ;
        RECT 131.690 197.095 132.010 197.155 ;
        RECT 133.545 197.110 133.835 197.155 ;
        RECT 134.080 197.155 137.055 197.295 ;
        RECT 123.870 196.955 124.190 197.015 ;
        RECT 134.080 196.955 134.220 197.155 ;
        RECT 136.765 197.110 137.055 197.155 ;
        RECT 137.225 197.110 137.515 197.340 ;
        RECT 139.065 197.110 139.355 197.340 ;
        RECT 139.510 197.295 139.830 197.355 ;
        RECT 140.905 197.295 141.195 197.340 ;
        RECT 139.510 197.155 141.195 197.295 ;
        RECT 121.660 196.815 124.190 196.955 ;
        RECT 119.730 196.755 120.050 196.815 ;
        RECT 121.125 196.770 121.415 196.815 ;
        RECT 123.870 196.755 124.190 196.815 ;
        RECT 124.420 196.815 134.220 196.955 ;
        RECT 136.290 196.955 136.610 197.015 ;
        RECT 137.300 196.955 137.440 197.110 ;
        RECT 139.140 196.955 139.280 197.110 ;
        RECT 139.510 197.095 139.830 197.155 ;
        RECT 140.905 197.110 141.195 197.155 ;
        RECT 142.730 197.095 143.050 197.355 ;
        RECT 144.660 197.340 144.800 197.835 ;
        RECT 144.585 197.110 144.875 197.340 ;
        RECT 136.290 196.815 137.440 196.955 ;
        RECT 137.760 196.815 139.280 196.955 ;
        RECT 76.965 196.475 80.400 196.615 ;
        RECT 76.965 196.430 77.255 196.475 ;
        RECT 81.550 196.415 81.870 196.675 ;
        RECT 91.225 196.615 91.515 196.660 ;
        RECT 92.590 196.615 92.910 196.675 ;
        RECT 91.225 196.475 92.910 196.615 ;
        RECT 93.140 196.615 93.280 196.755 ;
        RECT 124.420 196.675 124.560 196.815 ;
        RECT 136.290 196.755 136.610 196.815 ;
        RECT 99.950 196.615 100.270 196.675 ;
        RECT 93.140 196.475 100.270 196.615 ;
        RECT 91.225 196.430 91.515 196.475 ;
        RECT 92.590 196.415 92.910 196.475 ;
        RECT 99.950 196.415 100.270 196.475 ;
        RECT 100.410 196.615 100.730 196.675 ;
        RECT 105.010 196.615 105.330 196.675 ;
        RECT 100.410 196.475 105.330 196.615 ;
        RECT 100.410 196.415 100.730 196.475 ;
        RECT 105.010 196.415 105.330 196.475 ;
        RECT 105.470 196.415 105.790 196.675 ;
        RECT 106.390 196.415 106.710 196.675 ;
        RECT 110.545 196.615 110.835 196.660 ;
        RECT 111.910 196.615 112.230 196.675 ;
        RECT 110.545 196.475 112.230 196.615 ;
        RECT 110.545 196.430 110.835 196.475 ;
        RECT 111.910 196.415 112.230 196.475 ;
        RECT 113.750 196.615 114.070 196.675 ;
        RECT 121.585 196.615 121.875 196.660 ;
        RECT 113.750 196.475 121.875 196.615 ;
        RECT 113.750 196.415 114.070 196.475 ;
        RECT 121.585 196.430 121.875 196.475 ;
        RECT 124.330 196.415 124.650 196.675 ;
        RECT 127.090 196.615 127.410 196.675 ;
        RECT 127.565 196.615 127.855 196.660 ;
        RECT 127.090 196.475 127.855 196.615 ;
        RECT 127.090 196.415 127.410 196.475 ;
        RECT 127.565 196.430 127.855 196.475 ;
        RECT 128.010 196.615 128.330 196.675 ;
        RECT 128.485 196.615 128.775 196.660 ;
        RECT 128.010 196.475 128.775 196.615 ;
        RECT 128.010 196.415 128.330 196.475 ;
        RECT 128.485 196.430 128.775 196.475 ;
        RECT 131.690 196.415 132.010 196.675 ;
        RECT 132.150 196.615 132.470 196.675 ;
        RECT 135.845 196.615 136.135 196.660 ;
        RECT 132.150 196.475 136.135 196.615 ;
        RECT 132.150 196.415 132.470 196.475 ;
        RECT 135.845 196.430 136.135 196.475 ;
        RECT 137.210 196.615 137.530 196.675 ;
        RECT 137.760 196.615 137.900 196.815 ;
        RECT 137.210 196.475 137.900 196.615 ;
        RECT 137.210 196.415 137.530 196.475 ;
        RECT 138.130 196.415 138.450 196.675 ;
        RECT 139.050 196.615 139.370 196.675 ;
        RECT 139.985 196.615 140.275 196.660 ;
        RECT 139.050 196.475 140.275 196.615 ;
        RECT 139.050 196.415 139.370 196.475 ;
        RECT 139.985 196.430 140.275 196.475 ;
        RECT 141.810 196.415 142.130 196.675 ;
        RECT 143.650 196.415 143.970 196.675 ;
        RECT 13.860 195.795 147.720 196.275 ;
        RECT 14.850 195.595 15.170 195.655 ;
        RECT 17.625 195.595 17.915 195.640 ;
        RECT 29.585 195.595 29.875 195.640 ;
        RECT 14.850 195.455 17.915 195.595 ;
        RECT 14.850 195.395 15.170 195.455 ;
        RECT 17.625 195.410 17.915 195.455 ;
        RECT 20.460 195.455 29.875 195.595 ;
        RECT 20.460 195.300 20.600 195.455 ;
        RECT 29.585 195.410 29.875 195.455 ;
        RECT 30.950 195.595 31.270 195.655 ;
        RECT 35.565 195.595 35.855 195.640 ;
        RECT 36.010 195.595 36.330 195.655 ;
        RECT 30.950 195.455 35.320 195.595 ;
        RECT 30.950 195.395 31.270 195.455 ;
        RECT 20.385 195.070 20.675 195.300 ;
        RECT 22.665 195.255 23.315 195.300 ;
        RECT 26.265 195.255 26.555 195.300 ;
        RECT 22.665 195.115 26.555 195.255 ;
        RECT 22.665 195.070 23.315 195.115 ;
        RECT 25.965 195.070 26.555 195.115 ;
        RECT 28.650 195.255 28.970 195.315 ;
        RECT 30.030 195.255 30.350 195.315 ;
        RECT 31.425 195.255 31.715 195.300 ;
        RECT 34.630 195.255 34.950 195.315 ;
        RECT 28.650 195.115 34.950 195.255 ;
        RECT 25.965 194.975 26.255 195.070 ;
        RECT 28.650 195.055 28.970 195.115 ;
        RECT 30.030 195.055 30.350 195.115 ;
        RECT 31.425 195.070 31.715 195.115 ;
        RECT 34.630 195.055 34.950 195.115 ;
        RECT 35.180 195.255 35.320 195.455 ;
        RECT 35.565 195.455 36.330 195.595 ;
        RECT 35.565 195.410 35.855 195.455 ;
        RECT 36.010 195.395 36.330 195.455 ;
        RECT 36.945 195.595 37.235 195.640 ;
        RECT 38.770 195.595 39.090 195.655 ;
        RECT 36.945 195.455 39.090 195.595 ;
        RECT 36.945 195.410 37.235 195.455 ;
        RECT 38.770 195.395 39.090 195.455 ;
        RECT 43.370 195.595 43.690 195.655 ;
        RECT 46.145 195.595 46.435 195.640 ;
        RECT 43.370 195.455 46.435 195.595 ;
        RECT 43.370 195.395 43.690 195.455 ;
        RECT 46.145 195.410 46.435 195.455 ;
        RECT 48.430 195.595 48.750 195.655 ;
        RECT 49.825 195.595 50.115 195.640 ;
        RECT 48.430 195.455 50.115 195.595 ;
        RECT 48.430 195.395 48.750 195.455 ;
        RECT 49.825 195.410 50.115 195.455 ;
        RECT 51.650 195.395 51.970 195.655 ;
        RECT 52.110 195.395 52.430 195.655 ;
        RECT 54.870 195.595 55.190 195.655 ;
        RECT 53.120 195.455 55.190 195.595 ;
        RECT 37.850 195.255 38.170 195.315 ;
        RECT 35.180 195.115 38.170 195.255 ;
        RECT 16.690 194.715 17.010 194.975 ;
        RECT 18.070 194.915 18.390 194.975 ;
        RECT 18.545 194.915 18.835 194.960 ;
        RECT 18.070 194.775 18.835 194.915 ;
        RECT 18.070 194.715 18.390 194.775 ;
        RECT 18.545 194.730 18.835 194.775 ;
        RECT 18.990 194.715 19.310 194.975 ;
        RECT 19.470 194.915 19.760 194.960 ;
        RECT 21.305 194.915 21.595 194.960 ;
        RECT 24.885 194.915 25.175 194.960 ;
        RECT 19.470 194.775 25.175 194.915 ;
        RECT 19.470 194.730 19.760 194.775 ;
        RECT 21.305 194.730 21.595 194.775 ;
        RECT 24.885 194.730 25.175 194.775 ;
        RECT 25.890 194.755 26.255 194.975 ;
        RECT 29.570 194.915 29.890 194.975 ;
        RECT 30.505 194.915 30.795 194.960 ;
        RECT 29.570 194.775 30.795 194.915 ;
        RECT 25.890 194.715 26.210 194.755 ;
        RECT 29.570 194.715 29.890 194.775 ;
        RECT 30.505 194.730 30.795 194.775 ;
        RECT 30.950 194.715 31.270 194.975 ;
        RECT 32.345 194.915 32.635 194.960 ;
        RECT 32.805 194.915 33.095 194.960 ;
        RECT 33.710 194.915 34.030 194.975 ;
        RECT 32.345 194.775 34.030 194.915 ;
        RECT 32.345 194.730 32.635 194.775 ;
        RECT 32.805 194.730 33.095 194.775 ;
        RECT 29.125 194.575 29.415 194.620 ;
        RECT 32.420 194.575 32.560 194.730 ;
        RECT 33.710 194.715 34.030 194.775 ;
        RECT 34.185 194.915 34.475 194.960 ;
        RECT 35.180 194.915 35.320 195.115 ;
        RECT 37.850 195.055 38.170 195.115 ;
        RECT 34.185 194.775 35.320 194.915 ;
        RECT 35.550 194.915 35.870 194.975 ;
        RECT 36.485 194.915 36.775 194.960 ;
        RECT 36.930 194.915 37.250 194.975 ;
        RECT 38.860 194.960 39.000 195.395 ;
        RECT 41.530 195.255 41.850 195.315 ;
        RECT 50.270 195.255 50.590 195.315 ;
        RECT 39.320 195.115 44.520 195.255 ;
        RECT 39.320 194.960 39.460 195.115 ;
        RECT 41.530 195.055 41.850 195.115 ;
        RECT 35.550 194.775 37.250 194.915 ;
        RECT 34.185 194.730 34.475 194.775 ;
        RECT 35.550 194.715 35.870 194.775 ;
        RECT 36.485 194.730 36.775 194.775 ;
        RECT 36.930 194.715 37.250 194.775 ;
        RECT 38.785 194.730 39.075 194.960 ;
        RECT 39.245 194.730 39.535 194.960 ;
        RECT 29.125 194.435 32.560 194.575 ;
        RECT 38.860 194.575 39.000 194.730 ;
        RECT 40.610 194.715 40.930 194.975 ;
        RECT 41.070 194.915 41.390 194.975 ;
        RECT 44.380 194.960 44.520 195.115 ;
        RECT 46.680 195.115 50.590 195.255 ;
        RECT 46.680 194.960 46.820 195.115 ;
        RECT 50.270 195.055 50.590 195.115 ;
        RECT 42.925 194.915 43.215 194.960 ;
        RECT 41.070 194.775 43.215 194.915 ;
        RECT 41.070 194.715 41.390 194.775 ;
        RECT 42.925 194.730 43.215 194.775 ;
        RECT 44.305 194.730 44.595 194.960 ;
        RECT 46.605 194.730 46.895 194.960 ;
        RECT 47.510 194.715 47.830 194.975 ;
        RECT 52.110 194.915 52.430 194.975 ;
        RECT 53.120 194.960 53.260 195.455 ;
        RECT 54.870 195.395 55.190 195.455 ;
        RECT 55.790 195.595 56.110 195.655 ;
        RECT 55.790 195.455 58.780 195.595 ;
        RECT 55.790 195.395 56.110 195.455 ;
        RECT 56.250 195.255 56.570 195.315 ;
        RECT 54.500 195.115 56.570 195.255 ;
        RECT 53.045 194.915 53.335 194.960 ;
        RECT 52.110 194.775 53.335 194.915 ;
        RECT 52.110 194.715 52.430 194.775 ;
        RECT 53.045 194.730 53.335 194.775 ;
        RECT 53.490 194.715 53.810 194.975 ;
        RECT 54.500 194.960 54.640 195.115 ;
        RECT 56.250 195.055 56.570 195.115 ;
        RECT 56.725 195.255 57.015 195.300 ;
        RECT 58.090 195.255 58.410 195.315 ;
        RECT 56.725 195.115 58.410 195.255 ;
        RECT 56.725 195.070 57.015 195.115 ;
        RECT 58.090 195.055 58.410 195.115 ;
        RECT 54.425 194.730 54.715 194.960 ;
        RECT 55.330 194.715 55.650 194.975 ;
        RECT 58.640 194.960 58.780 195.455 ;
        RECT 59.010 195.395 59.330 195.655 ;
        RECT 59.470 195.595 59.790 195.655 ;
        RECT 59.470 195.455 60.160 195.595 ;
        RECT 59.470 195.395 59.790 195.455 ;
        RECT 59.100 195.255 59.240 195.395 ;
        RECT 60.020 195.300 60.160 195.455 ;
        RECT 61.310 195.395 61.630 195.655 ;
        RECT 62.230 195.595 62.550 195.655 ;
        RECT 80.630 195.595 80.950 195.655 ;
        RECT 85.230 195.595 85.550 195.655 ;
        RECT 87.990 195.595 88.310 195.655 ;
        RECT 110.990 195.595 111.310 195.655 ;
        RECT 62.230 195.455 80.950 195.595 ;
        RECT 62.230 195.395 62.550 195.455 ;
        RECT 80.630 195.395 80.950 195.455 ;
        RECT 81.640 195.455 88.310 195.595 ;
        RECT 59.945 195.255 60.235 195.300 ;
        RECT 67.305 195.255 67.595 195.300 ;
        RECT 68.210 195.255 68.530 195.315 ;
        RECT 59.100 195.115 59.700 195.255 ;
        RECT 57.185 194.730 57.475 194.960 ;
        RECT 58.565 194.915 58.855 194.960 ;
        RECT 59.010 194.915 59.330 194.975 ;
        RECT 59.560 194.960 59.700 195.115 ;
        RECT 59.945 195.115 66.140 195.255 ;
        RECT 59.945 195.070 60.235 195.115 ;
        RECT 58.565 194.775 59.330 194.915 ;
        RECT 58.565 194.730 58.855 194.775 ;
        RECT 43.370 194.575 43.690 194.635 ;
        RECT 44.765 194.575 45.055 194.620 ;
        RECT 38.860 194.435 43.140 194.575 ;
        RECT 29.125 194.390 29.415 194.435 ;
        RECT 14.390 194.235 14.710 194.295 ;
        RECT 15.785 194.235 16.075 194.280 ;
        RECT 14.390 194.095 16.075 194.235 ;
        RECT 14.390 194.035 14.710 194.095 ;
        RECT 15.785 194.050 16.075 194.095 ;
        RECT 19.875 194.235 20.165 194.280 ;
        RECT 21.765 194.235 22.055 194.280 ;
        RECT 24.885 194.235 25.175 194.280 ;
        RECT 19.875 194.095 25.175 194.235 ;
        RECT 19.875 194.050 20.165 194.095 ;
        RECT 21.765 194.050 22.055 194.095 ;
        RECT 24.885 194.050 25.175 194.095 ;
        RECT 25.430 194.235 25.750 194.295 ;
        RECT 25.430 194.095 35.780 194.235 ;
        RECT 25.430 194.035 25.750 194.095 ;
        RECT 27.730 193.895 28.050 193.955 ;
        RECT 33.250 193.895 33.570 193.955 ;
        RECT 27.730 193.755 33.570 193.895 ;
        RECT 35.640 193.895 35.780 194.095 ;
        RECT 39.230 194.035 39.550 194.295 ;
        RECT 43.000 194.235 43.140 194.435 ;
        RECT 43.370 194.435 45.055 194.575 ;
        RECT 43.370 194.375 43.690 194.435 ;
        RECT 44.765 194.390 45.055 194.435 ;
        RECT 47.970 194.575 48.290 194.635 ;
        RECT 48.445 194.575 48.735 194.620 ;
        RECT 47.970 194.435 48.735 194.575 ;
        RECT 47.970 194.375 48.290 194.435 ;
        RECT 48.445 194.390 48.735 194.435 ;
        RECT 49.365 194.390 49.655 194.620 ;
        RECT 52.570 194.575 52.890 194.635 ;
        RECT 53.965 194.575 54.255 194.620 ;
        RECT 55.420 194.575 55.560 194.715 ;
        RECT 52.570 194.435 54.255 194.575 ;
        RECT 49.440 194.235 49.580 194.390 ;
        RECT 52.570 194.375 52.890 194.435 ;
        RECT 53.965 194.390 54.255 194.435 ;
        RECT 54.560 194.435 55.560 194.575 ;
        RECT 57.260 194.575 57.400 194.730 ;
        RECT 59.010 194.715 59.330 194.775 ;
        RECT 59.485 194.730 59.775 194.960 ;
        RECT 59.560 194.575 59.700 194.730 ;
        RECT 60.390 194.715 60.710 194.975 ;
        RECT 66.000 194.960 66.140 195.115 ;
        RECT 67.305 195.115 68.530 195.255 ;
        RECT 67.305 195.070 67.595 195.115 ;
        RECT 68.210 195.055 68.530 195.115 ;
        RECT 68.670 195.255 68.990 195.315 ;
        RECT 72.805 195.255 73.455 195.300 ;
        RECT 76.405 195.255 76.695 195.300 ;
        RECT 68.670 195.115 76.695 195.255 ;
        RECT 68.670 195.055 68.990 195.115 ;
        RECT 72.805 195.070 73.455 195.115 ;
        RECT 76.105 195.070 76.695 195.115 ;
        RECT 76.950 195.255 77.270 195.315 ;
        RECT 79.265 195.255 79.555 195.300 ;
        RECT 81.090 195.255 81.410 195.315 ;
        RECT 76.950 195.115 81.410 195.255 ;
        RECT 65.925 194.915 66.215 194.960 ;
        RECT 65.925 194.775 66.600 194.915 ;
        RECT 65.925 194.730 66.215 194.775 ;
        RECT 65.450 194.575 65.770 194.635 ;
        RECT 57.260 194.435 59.240 194.575 ;
        RECT 59.560 194.435 65.770 194.575 ;
        RECT 54.560 194.235 54.700 194.435 ;
        RECT 43.000 194.095 44.980 194.235 ;
        RECT 49.440 194.095 54.700 194.235 ;
        RECT 54.870 194.235 55.190 194.295 ;
        RECT 57.260 194.235 57.400 194.435 ;
        RECT 54.870 194.095 57.400 194.235 ;
        RECT 40.610 193.895 40.930 193.955 ;
        RECT 44.840 193.940 44.980 194.095 ;
        RECT 54.870 194.035 55.190 194.095 ;
        RECT 35.640 193.755 40.930 193.895 ;
        RECT 27.730 193.695 28.050 193.755 ;
        RECT 33.250 193.695 33.570 193.755 ;
        RECT 40.610 193.695 40.930 193.755 ;
        RECT 44.765 193.710 45.055 193.940 ;
        RECT 47.050 193.695 47.370 193.955 ;
        RECT 53.490 193.895 53.810 193.955 ;
        RECT 55.790 193.895 56.110 193.955 ;
        RECT 53.490 193.755 56.110 193.895 ;
        RECT 53.490 193.695 53.810 193.755 ;
        RECT 55.790 193.695 56.110 193.755 ;
        RECT 58.090 193.695 58.410 193.955 ;
        RECT 59.100 193.895 59.240 194.435 ;
        RECT 65.450 194.375 65.770 194.435 ;
        RECT 59.470 194.235 59.790 194.295 ;
        RECT 63.150 194.235 63.470 194.295 ;
        RECT 59.470 194.095 63.470 194.235 ;
        RECT 59.470 194.035 59.790 194.095 ;
        RECT 63.150 194.035 63.470 194.095 ;
        RECT 62.230 193.895 62.550 193.955 ;
        RECT 59.100 193.755 62.550 193.895 ;
        RECT 66.460 193.895 66.600 194.775 ;
        RECT 66.830 194.715 67.150 194.975 ;
        RECT 67.750 194.715 68.070 194.975 ;
        RECT 69.130 194.715 69.450 194.975 ;
        RECT 69.610 194.915 69.900 194.960 ;
        RECT 71.445 194.915 71.735 194.960 ;
        RECT 75.025 194.915 75.315 194.960 ;
        RECT 69.610 194.775 75.315 194.915 ;
        RECT 69.610 194.730 69.900 194.775 ;
        RECT 71.445 194.730 71.735 194.775 ;
        RECT 75.025 194.730 75.315 194.775 ;
        RECT 76.105 194.755 76.395 195.070 ;
        RECT 76.950 195.055 77.270 195.115 ;
        RECT 79.265 195.070 79.555 195.115 ;
        RECT 81.090 195.055 81.410 195.115 ;
        RECT 80.170 194.915 80.490 194.975 ;
        RECT 81.640 194.915 81.780 195.455 ;
        RECT 85.230 195.395 85.550 195.455 ;
        RECT 87.990 195.395 88.310 195.455 ;
        RECT 91.760 195.455 111.310 195.595 ;
        RECT 82.010 195.255 82.330 195.315 ;
        RECT 82.585 195.255 82.875 195.300 ;
        RECT 85.825 195.255 86.475 195.300 ;
        RECT 82.010 195.115 86.475 195.255 ;
        RECT 82.010 195.055 82.330 195.115 ;
        RECT 82.585 195.070 83.175 195.115 ;
        RECT 85.825 195.070 86.475 195.115 ;
        RECT 80.170 194.775 81.780 194.915 ;
        RECT 80.170 194.715 80.490 194.775 ;
        RECT 82.885 194.755 83.175 195.070 ;
        RECT 91.760 194.960 91.900 195.455 ;
        RECT 110.990 195.395 111.310 195.455 ;
        RECT 112.370 195.595 112.690 195.655 ;
        RECT 113.305 195.595 113.595 195.640 ;
        RECT 112.370 195.455 113.595 195.595 ;
        RECT 112.370 195.395 112.690 195.455 ;
        RECT 113.305 195.410 113.595 195.455 ;
        RECT 115.590 195.595 115.910 195.655 ;
        RECT 117.445 195.595 117.735 195.640 ;
        RECT 115.590 195.455 117.735 195.595 ;
        RECT 115.590 195.395 115.910 195.455 ;
        RECT 117.445 195.410 117.735 195.455 ;
        RECT 126.170 195.595 126.490 195.655 ;
        RECT 128.930 195.595 129.250 195.655 ;
        RECT 133.990 195.595 134.310 195.655 ;
        RECT 126.170 195.455 129.250 195.595 ;
        RECT 126.170 195.395 126.490 195.455 ;
        RECT 128.930 195.395 129.250 195.455 ;
        RECT 129.480 195.455 134.310 195.595 ;
        RECT 95.345 195.255 95.995 195.300 ;
        RECT 98.945 195.255 99.235 195.300 ;
        RECT 95.345 195.115 99.235 195.255 ;
        RECT 95.345 195.070 95.995 195.115 ;
        RECT 98.645 195.070 99.235 195.115 ;
        RECT 99.490 195.255 99.810 195.315 ;
        RECT 111.080 195.255 111.220 195.395 ;
        RECT 116.510 195.255 116.830 195.315 ;
        RECT 122.030 195.255 122.350 195.315 ;
        RECT 99.490 195.115 104.780 195.255 ;
        RECT 111.080 195.115 122.350 195.255 ;
        RECT 98.645 194.975 98.935 195.070 ;
        RECT 99.490 195.055 99.810 195.115 ;
        RECT 104.640 194.975 104.780 195.115 ;
        RECT 116.510 195.055 116.830 195.115 ;
        RECT 83.965 194.915 84.255 194.960 ;
        RECT 87.545 194.915 87.835 194.960 ;
        RECT 89.380 194.915 89.670 194.960 ;
        RECT 83.965 194.775 89.670 194.915 ;
        RECT 83.965 194.730 84.255 194.775 ;
        RECT 87.545 194.730 87.835 194.775 ;
        RECT 89.380 194.730 89.670 194.775 ;
        RECT 89.845 194.915 90.135 194.960 ;
        RECT 91.685 194.915 91.975 194.960 ;
        RECT 89.845 194.775 91.975 194.915 ;
        RECT 89.845 194.730 90.135 194.775 ;
        RECT 91.685 194.730 91.975 194.775 ;
        RECT 92.150 194.915 92.440 194.960 ;
        RECT 93.985 194.915 94.275 194.960 ;
        RECT 97.565 194.915 97.855 194.960 ;
        RECT 92.150 194.775 97.855 194.915 ;
        RECT 92.150 194.730 92.440 194.775 ;
        RECT 93.985 194.730 94.275 194.775 ;
        RECT 97.565 194.730 97.855 194.775 ;
        RECT 98.570 194.755 98.935 194.975 ;
        RECT 103.185 194.915 103.475 194.960 ;
        RECT 99.120 194.775 103.475 194.915 ;
        RECT 98.570 194.715 98.890 194.755 ;
        RECT 70.525 194.575 70.815 194.620 ;
        RECT 68.760 194.435 70.815 194.575 ;
        RECT 68.760 194.280 68.900 194.435 ;
        RECT 70.525 194.390 70.815 194.435 ;
        RECT 74.190 194.575 74.510 194.635 ;
        RECT 78.790 194.575 79.110 194.635 ;
        RECT 79.725 194.575 80.015 194.620 ;
        RECT 74.190 194.435 80.015 194.575 ;
        RECT 74.190 194.375 74.510 194.435 ;
        RECT 78.790 194.375 79.110 194.435 ;
        RECT 79.725 194.390 80.015 194.435 ;
        RECT 84.770 194.575 85.090 194.635 ;
        RECT 88.465 194.575 88.755 194.620 ;
        RECT 84.770 194.435 88.755 194.575 ;
        RECT 84.770 194.375 85.090 194.435 ;
        RECT 88.465 194.390 88.755 194.435 ;
        RECT 93.050 194.375 93.370 194.635 ;
        RECT 96.730 194.575 97.050 194.635 ;
        RECT 99.120 194.575 99.260 194.775 ;
        RECT 103.185 194.730 103.475 194.775 ;
        RECT 103.630 194.715 103.950 194.975 ;
        RECT 104.550 194.715 104.870 194.975 ;
        RECT 105.930 194.915 106.250 194.975 ;
        RECT 106.865 194.915 107.155 194.960 ;
        RECT 105.930 194.775 107.155 194.915 ;
        RECT 105.930 194.715 106.250 194.775 ;
        RECT 106.865 194.730 107.155 194.775 ;
        RECT 109.150 194.715 109.470 194.975 ;
        RECT 110.530 194.915 110.850 194.975 ;
        RECT 111.005 194.915 111.295 194.960 ;
        RECT 110.530 194.775 111.295 194.915 ;
        RECT 110.530 194.715 110.850 194.775 ;
        RECT 111.005 194.730 111.295 194.775 ;
        RECT 96.730 194.435 99.260 194.575 ;
        RECT 99.950 194.575 100.270 194.635 ;
        RECT 101.805 194.575 102.095 194.620 ;
        RECT 103.720 194.575 103.860 194.715 ;
        RECT 99.950 194.435 102.095 194.575 ;
        RECT 96.730 194.375 97.050 194.435 ;
        RECT 99.950 194.375 100.270 194.435 ;
        RECT 101.805 194.390 102.095 194.435 ;
        RECT 102.340 194.435 103.860 194.575 ;
        RECT 105.470 194.575 105.790 194.635 ;
        RECT 107.325 194.575 107.615 194.620 ;
        RECT 105.470 194.435 107.615 194.575 ;
        RECT 68.685 194.050 68.975 194.280 ;
        RECT 70.015 194.235 70.305 194.280 ;
        RECT 71.905 194.235 72.195 194.280 ;
        RECT 75.025 194.235 75.315 194.280 ;
        RECT 70.015 194.095 75.315 194.235 ;
        RECT 70.015 194.050 70.305 194.095 ;
        RECT 71.905 194.050 72.195 194.095 ;
        RECT 75.025 194.050 75.315 194.095 ;
        RECT 83.965 194.235 84.255 194.280 ;
        RECT 87.085 194.235 87.375 194.280 ;
        RECT 88.975 194.235 89.265 194.280 ;
        RECT 83.965 194.095 89.265 194.235 ;
        RECT 83.965 194.050 84.255 194.095 ;
        RECT 87.085 194.050 87.375 194.095 ;
        RECT 88.975 194.050 89.265 194.095 ;
        RECT 92.555 194.235 92.845 194.280 ;
        RECT 94.445 194.235 94.735 194.280 ;
        RECT 97.565 194.235 97.855 194.280 ;
        RECT 92.555 194.095 97.855 194.235 ;
        RECT 92.555 194.050 92.845 194.095 ;
        RECT 94.445 194.050 94.735 194.095 ;
        RECT 97.565 194.050 97.855 194.095 ;
        RECT 98.570 194.235 98.890 194.295 ;
        RECT 100.410 194.235 100.730 194.295 ;
        RECT 102.340 194.235 102.480 194.435 ;
        RECT 105.470 194.375 105.790 194.435 ;
        RECT 107.325 194.390 107.615 194.435 ;
        RECT 109.610 194.375 109.930 194.635 ;
        RECT 111.080 194.575 111.220 194.730 ;
        RECT 111.450 194.715 111.770 194.975 ;
        RECT 112.370 194.715 112.690 194.975 ;
        RECT 113.750 194.715 114.070 194.975 ;
        RECT 114.685 194.915 114.975 194.960 ;
        RECT 114.300 194.775 114.975 194.915 ;
        RECT 114.300 194.575 114.440 194.775 ;
        RECT 114.685 194.730 114.975 194.775 ;
        RECT 115.145 194.730 115.435 194.960 ;
        RECT 111.080 194.435 114.440 194.575 ;
        RECT 115.220 194.575 115.360 194.730 ;
        RECT 115.590 194.715 115.910 194.975 ;
        RECT 119.730 194.915 120.050 194.975 ;
        RECT 120.280 194.960 120.420 195.115 ;
        RECT 122.030 195.055 122.350 195.115 ;
        RECT 123.865 195.255 124.515 195.300 ;
        RECT 127.465 195.255 127.755 195.300 ;
        RECT 123.865 195.115 127.755 195.255 ;
        RECT 123.865 195.070 124.515 195.115 ;
        RECT 127.165 195.070 127.755 195.115 ;
        RECT 117.980 194.775 120.050 194.915 ;
        RECT 117.980 194.575 118.120 194.775 ;
        RECT 119.730 194.715 120.050 194.775 ;
        RECT 120.205 194.730 120.495 194.960 ;
        RECT 120.670 194.915 120.960 194.960 ;
        RECT 122.505 194.915 122.795 194.960 ;
        RECT 126.085 194.915 126.375 194.960 ;
        RECT 120.670 194.775 126.375 194.915 ;
        RECT 120.670 194.730 120.960 194.775 ;
        RECT 122.505 194.730 122.795 194.775 ;
        RECT 126.085 194.730 126.375 194.775 ;
        RECT 126.630 194.915 126.950 194.975 ;
        RECT 127.165 194.915 127.455 195.070 ;
        RECT 126.630 194.775 127.455 194.915 ;
        RECT 126.630 194.715 126.950 194.775 ;
        RECT 127.165 194.755 127.455 194.775 ;
        RECT 115.220 194.435 118.120 194.575 ;
        RECT 98.570 194.095 100.730 194.235 ;
        RECT 98.570 194.035 98.890 194.095 ;
        RECT 100.410 194.035 100.730 194.095 ;
        RECT 100.960 194.095 102.480 194.235 ;
        RECT 102.710 194.235 103.030 194.295 ;
        RECT 105.945 194.235 106.235 194.280 ;
        RECT 115.220 194.235 115.360 194.435 ;
        RECT 118.350 194.375 118.670 194.635 ;
        RECT 118.810 194.375 119.130 194.635 ;
        RECT 119.270 194.375 119.590 194.635 ;
        RECT 121.585 194.575 121.875 194.620 ;
        RECT 120.280 194.435 121.875 194.575 ;
        RECT 102.710 194.095 106.235 194.235 ;
        RECT 70.510 193.895 70.830 193.955 ;
        RECT 66.460 193.755 70.830 193.895 ;
        RECT 62.230 193.695 62.550 193.755 ;
        RECT 70.510 193.695 70.830 193.755 ;
        RECT 72.350 193.895 72.670 193.955 ;
        RECT 82.930 193.895 83.250 193.955 ;
        RECT 91.670 193.895 91.990 193.955 ;
        RECT 100.960 193.895 101.100 194.095 ;
        RECT 102.710 194.035 103.030 194.095 ;
        RECT 105.945 194.050 106.235 194.095 ;
        RECT 111.540 194.095 115.360 194.235 ;
        RECT 116.525 194.235 116.815 194.280 ;
        RECT 120.280 194.235 120.420 194.435 ;
        RECT 121.585 194.390 121.875 194.435 ;
        RECT 123.870 194.575 124.190 194.635 ;
        RECT 127.180 194.575 127.320 194.755 ;
        RECT 129.480 194.575 129.620 195.455 ;
        RECT 133.990 195.395 134.310 195.455 ;
        RECT 134.450 195.595 134.770 195.655 ;
        RECT 136.765 195.595 137.055 195.640 ;
        RECT 134.450 195.455 137.055 195.595 ;
        RECT 134.450 195.395 134.770 195.455 ;
        RECT 136.765 195.410 137.055 195.455 ;
        RECT 145.490 195.395 145.810 195.655 ;
        RECT 132.610 195.055 132.930 195.315 ;
        RECT 130.785 194.730 131.075 194.960 ;
        RECT 131.230 194.915 131.550 194.975 ;
        RECT 131.705 194.915 131.995 194.960 ;
        RECT 131.230 194.775 131.995 194.915 ;
        RECT 123.870 194.435 129.620 194.575 ;
        RECT 130.860 194.575 131.000 194.730 ;
        RECT 131.230 194.715 131.550 194.775 ;
        RECT 131.705 194.730 131.995 194.775 ;
        RECT 132.165 194.915 132.455 194.960 ;
        RECT 132.700 194.915 132.840 195.055 ;
        RECT 132.165 194.775 132.840 194.915 ;
        RECT 132.165 194.730 132.455 194.775 ;
        RECT 133.070 194.715 133.390 194.975 ;
        RECT 133.530 194.715 133.850 194.975 ;
        RECT 134.005 194.730 134.295 194.960 ;
        RECT 132.610 194.575 132.930 194.635 ;
        RECT 130.860 194.435 132.930 194.575 ;
        RECT 133.160 194.575 133.300 194.715 ;
        RECT 134.080 194.575 134.220 194.730 ;
        RECT 134.910 194.715 135.230 194.975 ;
        RECT 136.750 194.915 137.070 194.975 ;
        RECT 137.685 194.915 137.975 194.960 ;
        RECT 136.750 194.775 137.975 194.915 ;
        RECT 136.750 194.715 137.070 194.775 ;
        RECT 137.685 194.730 137.975 194.775 ;
        RECT 138.145 194.730 138.435 194.960 ;
        RECT 133.160 194.435 134.220 194.575 ;
        RECT 135.845 194.575 136.135 194.620 ;
        RECT 138.220 194.575 138.360 194.730 ;
        RECT 140.890 194.715 141.210 194.975 ;
        RECT 143.190 194.715 143.510 194.975 ;
        RECT 144.125 194.730 144.415 194.960 ;
        RECT 135.845 194.435 138.360 194.575 ;
        RECT 140.430 194.575 140.750 194.635 ;
        RECT 143.650 194.575 143.970 194.635 ;
        RECT 144.200 194.575 144.340 194.730 ;
        RECT 144.570 194.715 144.890 194.975 ;
        RECT 140.430 194.435 144.340 194.575 ;
        RECT 123.870 194.375 124.190 194.435 ;
        RECT 132.610 194.375 132.930 194.435 ;
        RECT 135.845 194.390 136.135 194.435 ;
        RECT 140.430 194.375 140.750 194.435 ;
        RECT 143.650 194.375 143.970 194.435 ;
        RECT 116.525 194.095 120.420 194.235 ;
        RECT 121.075 194.235 121.365 194.280 ;
        RECT 122.965 194.235 123.255 194.280 ;
        RECT 126.085 194.235 126.375 194.280 ;
        RECT 121.075 194.095 126.375 194.235 ;
        RECT 111.540 193.955 111.680 194.095 ;
        RECT 116.525 194.050 116.815 194.095 ;
        RECT 121.075 194.050 121.365 194.095 ;
        RECT 122.965 194.050 123.255 194.095 ;
        RECT 126.085 194.050 126.375 194.095 ;
        RECT 128.930 194.235 129.250 194.295 ;
        RECT 130.310 194.235 130.630 194.295 ;
        RECT 131.245 194.235 131.535 194.280 ;
        RECT 128.930 194.095 131.535 194.235 ;
        RECT 128.930 194.035 129.250 194.095 ;
        RECT 130.310 194.035 130.630 194.095 ;
        RECT 131.245 194.050 131.535 194.095 ;
        RECT 133.530 194.235 133.850 194.295 ;
        RECT 139.065 194.235 139.355 194.280 ;
        RECT 143.205 194.235 143.495 194.280 ;
        RECT 133.530 194.095 139.355 194.235 ;
        RECT 72.350 193.755 101.100 193.895 ;
        RECT 72.350 193.695 72.670 193.755 ;
        RECT 82.930 193.695 83.250 193.755 ;
        RECT 91.670 193.695 91.990 193.755 ;
        RECT 102.250 193.695 102.570 193.955 ;
        RECT 103.170 193.895 103.490 193.955 ;
        RECT 103.645 193.895 103.935 193.940 ;
        RECT 103.170 193.755 103.935 193.895 ;
        RECT 103.170 193.695 103.490 193.755 ;
        RECT 103.645 193.710 103.935 193.755 ;
        RECT 104.090 193.895 104.410 193.955 ;
        RECT 111.450 193.895 111.770 193.955 ;
        RECT 104.090 193.755 111.770 193.895 ;
        RECT 104.090 193.695 104.410 193.755 ;
        RECT 111.450 193.695 111.770 193.755 ;
        RECT 117.890 193.895 118.210 193.955 ;
        RECT 129.865 193.895 130.155 193.940 ;
        RECT 117.890 193.755 130.155 193.895 ;
        RECT 131.320 193.895 131.460 194.050 ;
        RECT 133.530 194.035 133.850 194.095 ;
        RECT 139.065 194.050 139.355 194.095 ;
        RECT 139.600 194.095 143.495 194.235 ;
        RECT 139.600 193.895 139.740 194.095 ;
        RECT 143.205 194.050 143.495 194.095 ;
        RECT 131.320 193.755 139.740 193.895 ;
        RECT 141.825 193.895 142.115 193.940 ;
        RECT 142.730 193.895 143.050 193.955 ;
        RECT 141.825 193.755 143.050 193.895 ;
        RECT 117.890 193.695 118.210 193.755 ;
        RECT 129.865 193.710 130.155 193.755 ;
        RECT 141.825 193.710 142.115 193.755 ;
        RECT 142.730 193.695 143.050 193.755 ;
        RECT 13.860 193.075 147.720 193.555 ;
        RECT 15.770 192.675 16.090 192.935 ;
        RECT 17.610 192.675 17.930 192.935 ;
        RECT 22.070 192.735 26.120 192.875 ;
        RECT 14.850 192.535 15.170 192.595 ;
        RECT 21.305 192.535 21.595 192.580 ;
        RECT 14.850 192.395 21.595 192.535 ;
        RECT 14.850 192.335 15.170 192.395 ;
        RECT 21.305 192.350 21.595 192.395 ;
        RECT 13.930 192.195 14.250 192.255 ;
        RECT 22.070 192.195 22.210 192.735 ;
        RECT 25.980 192.535 26.120 192.735 ;
        RECT 27.270 192.675 27.590 192.935 ;
        RECT 36.025 192.690 36.315 192.920 ;
        RECT 36.945 192.875 37.235 192.920 ;
        RECT 37.390 192.875 37.710 192.935 ;
        RECT 36.945 192.735 37.710 192.875 ;
        RECT 36.945 192.690 37.235 192.735 ;
        RECT 32.805 192.535 33.095 192.580 ;
        RECT 25.980 192.395 33.095 192.535 ;
        RECT 36.100 192.535 36.240 192.690 ;
        RECT 37.390 192.675 37.710 192.735 ;
        RECT 37.865 192.875 38.155 192.920 ;
        RECT 38.310 192.875 38.630 192.935 ;
        RECT 37.865 192.735 38.630 192.875 ;
        RECT 37.865 192.690 38.155 192.735 ;
        RECT 38.310 192.675 38.630 192.735 ;
        RECT 41.530 192.875 41.850 192.935 ;
        RECT 42.465 192.875 42.755 192.920 ;
        RECT 41.530 192.735 42.755 192.875 ;
        RECT 41.530 192.675 41.850 192.735 ;
        RECT 42.465 192.690 42.755 192.735 ;
        RECT 43.920 192.735 55.100 192.875 ;
        RECT 40.165 192.535 40.455 192.580 ;
        RECT 36.100 192.395 40.455 192.535 ;
        RECT 32.805 192.350 33.095 192.395 ;
        RECT 40.165 192.350 40.455 192.395 ;
        RECT 40.610 192.535 40.930 192.595 ;
        RECT 43.920 192.535 44.060 192.735 ;
        RECT 40.610 192.395 44.060 192.535 ;
        RECT 40.610 192.335 40.930 192.395 ;
        RECT 32.330 192.195 32.650 192.255 ;
        RECT 13.930 192.055 22.210 192.195 ;
        RECT 24.600 192.055 32.650 192.195 ;
        RECT 13.930 191.995 14.250 192.055 ;
        RECT 16.690 191.655 17.010 191.915 ;
        RECT 18.545 191.855 18.835 191.900 ;
        RECT 19.910 191.855 20.230 191.915 ;
        RECT 18.545 191.715 20.230 191.855 ;
        RECT 18.545 191.670 18.835 191.715 ;
        RECT 19.910 191.655 20.230 191.715 ;
        RECT 20.370 191.655 20.690 191.915 ;
        RECT 22.225 191.855 22.515 191.900 ;
        RECT 24.600 191.855 24.740 192.055 ;
        RECT 32.330 191.995 32.650 192.055 ;
        RECT 33.250 192.195 33.570 192.255 ;
        RECT 35.565 192.195 35.855 192.240 ;
        RECT 37.850 192.195 38.170 192.255 ;
        RECT 43.370 192.195 43.690 192.255 ;
        RECT 33.250 192.055 34.400 192.195 ;
        RECT 33.250 191.995 33.570 192.055 ;
        RECT 22.225 191.715 24.740 191.855 ;
        RECT 22.225 191.670 22.515 191.715 ;
        RECT 24.970 191.655 25.290 191.915 ;
        RECT 28.205 191.670 28.495 191.900 ;
        RECT 23.130 191.515 23.450 191.575 ;
        RECT 23.605 191.515 23.895 191.560 ;
        RECT 23.130 191.375 23.895 191.515 ;
        RECT 23.130 191.315 23.450 191.375 ;
        RECT 23.605 191.330 23.895 191.375 ;
        RECT 24.525 191.515 24.815 191.560 ;
        RECT 26.810 191.515 27.130 191.575 ;
        RECT 24.525 191.375 27.130 191.515 ;
        RECT 28.280 191.515 28.420 191.670 ;
        RECT 28.650 191.655 28.970 191.915 ;
        RECT 29.110 191.655 29.430 191.915 ;
        RECT 30.045 191.855 30.335 191.900 ;
        RECT 31.410 191.855 31.730 191.915 ;
        RECT 30.045 191.715 31.730 191.855 ;
        RECT 30.045 191.670 30.335 191.715 ;
        RECT 31.410 191.655 31.730 191.715 ;
        RECT 31.870 191.655 32.190 191.915 ;
        RECT 32.790 191.655 33.110 191.915 ;
        RECT 33.710 191.655 34.030 191.915 ;
        RECT 34.260 191.900 34.400 192.055 ;
        RECT 35.565 192.055 43.690 192.195 ;
        RECT 35.565 192.010 35.855 192.055 ;
        RECT 37.850 191.995 38.170 192.055 ;
        RECT 43.370 191.995 43.690 192.055 ;
        RECT 34.185 191.670 34.475 191.900 ;
        RECT 38.770 191.655 39.090 191.915 ;
        RECT 41.085 191.670 41.375 191.900 ;
        RECT 32.880 191.515 33.020 191.655 ;
        RECT 28.280 191.375 33.020 191.515 ;
        RECT 34.630 191.515 34.950 191.575 ;
        RECT 41.160 191.515 41.300 191.670 ;
        RECT 41.530 191.655 41.850 191.915 ;
        RECT 43.920 191.900 44.060 192.395 ;
        RECT 48.445 192.535 48.735 192.580 ;
        RECT 49.810 192.535 50.130 192.595 ;
        RECT 53.030 192.535 53.350 192.595 ;
        RECT 48.445 192.395 50.130 192.535 ;
        RECT 48.445 192.350 48.735 192.395 ;
        RECT 49.810 192.335 50.130 192.395 ;
        RECT 51.280 192.395 53.350 192.535 ;
        RECT 47.525 192.195 47.815 192.240 ;
        RECT 51.280 192.195 51.420 192.395 ;
        RECT 53.030 192.335 53.350 192.395 ;
        RECT 47.525 192.055 51.420 192.195 ;
        RECT 54.960 192.195 55.100 192.735 ;
        RECT 55.790 192.675 56.110 192.935 ;
        RECT 70.525 192.875 70.815 192.920 ;
        RECT 70.970 192.875 71.290 192.935 ;
        RECT 56.800 192.735 62.000 192.875 ;
        RECT 56.800 192.195 56.940 192.735 ;
        RECT 54.960 192.055 56.940 192.195 ;
        RECT 47.525 192.010 47.815 192.055 ;
        RECT 42.925 191.670 43.215 191.900 ;
        RECT 43.845 191.670 44.135 191.900 ;
        RECT 44.305 191.670 44.595 191.900 ;
        RECT 46.605 191.670 46.895 191.900 ;
        RECT 47.065 191.670 47.355 191.900 ;
        RECT 48.430 191.855 48.750 191.915 ;
        RECT 48.905 191.855 49.195 191.900 ;
        RECT 48.430 191.715 49.195 191.855 ;
        RECT 34.630 191.375 41.300 191.515 ;
        RECT 24.525 191.330 24.815 191.375 ;
        RECT 26.810 191.315 27.130 191.375 ;
        RECT 34.630 191.315 34.950 191.375 ;
        RECT 13.470 191.175 13.790 191.235 ;
        RECT 19.465 191.175 19.755 191.220 ;
        RECT 13.470 191.035 19.755 191.175 ;
        RECT 13.470 190.975 13.790 191.035 ;
        RECT 19.465 190.990 19.755 191.035 ;
        RECT 25.905 191.175 26.195 191.220 ;
        RECT 27.730 191.175 28.050 191.235 ;
        RECT 25.905 191.035 28.050 191.175 ;
        RECT 25.905 190.990 26.195 191.035 ;
        RECT 27.730 190.975 28.050 191.035 ;
        RECT 28.190 191.175 28.510 191.235 ;
        RECT 30.965 191.175 31.255 191.220 ;
        RECT 28.190 191.035 31.255 191.175 ;
        RECT 28.190 190.975 28.510 191.035 ;
        RECT 30.965 190.990 31.255 191.035 ;
        RECT 31.410 191.175 31.730 191.235 ;
        RECT 43.000 191.175 43.140 191.670 ;
        RECT 43.385 191.515 43.675 191.560 ;
        RECT 44.380 191.515 44.520 191.670 ;
        RECT 46.680 191.515 46.820 191.670 ;
        RECT 43.385 191.375 44.520 191.515 ;
        RECT 44.840 191.375 46.820 191.515 ;
        RECT 47.140 191.515 47.280 191.670 ;
        RECT 48.430 191.655 48.750 191.715 ;
        RECT 48.905 191.670 49.195 191.715 ;
        RECT 49.810 191.655 50.130 191.915 ;
        RECT 50.745 191.855 51.035 191.900 ;
        RECT 52.110 191.855 52.430 191.915 ;
        RECT 54.960 191.900 55.100 192.055 ;
        RECT 57.170 191.995 57.490 192.255 ;
        RECT 57.735 192.195 58.025 192.240 ;
        RECT 57.720 192.085 58.025 192.195 ;
        RECT 57.630 192.010 58.025 192.085 ;
        RECT 61.860 192.195 62.000 192.735 ;
        RECT 70.525 192.735 71.290 192.875 ;
        RECT 70.525 192.690 70.815 192.735 ;
        RECT 70.970 192.675 71.290 192.735 ;
        RECT 75.110 192.875 75.430 192.935 ;
        RECT 75.585 192.875 75.875 192.920 ;
        RECT 79.710 192.875 80.030 192.935 ;
        RECT 75.110 192.735 80.030 192.875 ;
        RECT 75.110 192.675 75.430 192.735 ;
        RECT 75.585 192.690 75.875 192.735 ;
        RECT 79.710 192.675 80.030 192.735 ;
        RECT 81.565 192.875 81.855 192.920 ;
        RECT 84.770 192.875 85.090 192.935 ;
        RECT 81.565 192.735 85.090 192.875 ;
        RECT 81.565 192.690 81.855 192.735 ;
        RECT 84.770 192.675 85.090 192.735 ;
        RECT 86.150 192.675 86.470 192.935 ;
        RECT 90.305 192.875 90.595 192.920 ;
        RECT 93.050 192.875 93.370 192.935 ;
        RECT 90.305 192.735 93.370 192.875 ;
        RECT 90.305 192.690 90.595 192.735 ;
        RECT 93.050 192.675 93.370 192.735 ;
        RECT 97.190 192.675 97.510 192.935 ;
        RECT 110.070 192.875 110.390 192.935 ;
        RECT 104.870 192.735 110.390 192.875 ;
        RECT 73.285 192.535 73.575 192.580 ;
        RECT 73.285 192.395 76.720 192.535 ;
        RECT 73.285 192.350 73.575 192.395 ;
        RECT 76.580 192.240 76.720 192.395 ;
        RECT 76.950 192.335 77.270 192.595 ;
        RECT 83.850 192.535 84.170 192.595 ;
        RECT 94.430 192.535 94.750 192.595 ;
        RECT 97.650 192.535 97.970 192.595 ;
        RECT 104.870 192.535 105.010 192.735 ;
        RECT 110.070 192.675 110.390 192.735 ;
        RECT 110.530 192.875 110.850 192.935 ;
        RECT 115.605 192.875 115.895 192.920 ;
        RECT 110.530 192.735 115.895 192.875 ;
        RECT 110.530 192.675 110.850 192.735 ;
        RECT 115.605 192.690 115.895 192.735 ;
        RECT 118.350 192.675 118.670 192.935 ;
        RECT 119.730 192.875 120.050 192.935 ;
        RECT 126.645 192.875 126.935 192.920 ;
        RECT 119.730 192.735 126.935 192.875 ;
        RECT 119.730 192.675 120.050 192.735 ;
        RECT 126.645 192.690 126.935 192.735 ;
        RECT 128.945 192.875 129.235 192.920 ;
        RECT 138.130 192.875 138.450 192.935 ;
        RECT 128.945 192.735 138.450 192.875 ;
        RECT 128.945 192.690 129.235 192.735 ;
        RECT 138.130 192.675 138.450 192.735 ;
        RECT 140.890 192.675 141.210 192.935 ;
        RECT 82.100 192.395 84.170 192.535 ;
        RECT 71.445 192.195 71.735 192.240 ;
        RECT 61.860 192.055 68.900 192.195 ;
        RECT 50.745 191.715 52.430 191.855 ;
        RECT 50.745 191.670 51.035 191.715 ;
        RECT 52.110 191.655 52.430 191.715 ;
        RECT 53.965 191.670 54.255 191.900 ;
        RECT 54.885 191.670 55.175 191.900 ;
        RECT 55.790 191.855 56.110 191.915 ;
        RECT 56.760 191.855 57.050 191.900 ;
        RECT 55.790 191.715 57.050 191.855 ;
        RECT 57.630 191.825 57.950 192.010 ;
        RECT 50.285 191.515 50.575 191.560 ;
        RECT 52.570 191.515 52.890 191.575 ;
        RECT 47.140 191.375 52.890 191.515 ;
        RECT 54.040 191.515 54.180 191.670 ;
        RECT 55.790 191.655 56.110 191.715 ;
        RECT 56.760 191.670 57.050 191.715 ;
        RECT 58.550 191.655 58.870 191.915 ;
        RECT 59.930 191.855 60.250 191.915 ;
        RECT 61.860 191.900 62.000 192.055 ;
        RECT 61.325 191.855 61.615 191.900 ;
        RECT 59.930 191.715 61.615 191.855 ;
        RECT 59.930 191.655 60.250 191.715 ;
        RECT 61.325 191.670 61.615 191.715 ;
        RECT 61.785 191.670 62.075 191.900 ;
        RECT 62.690 191.655 63.010 191.915 ;
        RECT 63.150 191.655 63.470 191.915 ;
        RECT 64.160 191.900 64.300 192.055 ;
        RECT 64.085 191.670 64.375 191.900 ;
        RECT 65.925 191.670 66.215 191.900 ;
        RECT 56.250 191.515 56.570 191.575 ;
        RECT 54.040 191.375 56.570 191.515 ;
        RECT 43.385 191.330 43.675 191.375 ;
        RECT 44.840 191.175 44.980 191.375 ;
        RECT 31.410 191.035 44.980 191.175 ;
        RECT 45.225 191.175 45.515 191.220 ;
        RECT 46.130 191.175 46.450 191.235 ;
        RECT 45.225 191.035 46.450 191.175 ;
        RECT 46.680 191.175 46.820 191.375 ;
        RECT 50.285 191.330 50.575 191.375 ;
        RECT 52.570 191.315 52.890 191.375 ;
        RECT 56.250 191.315 56.570 191.375 ;
        RECT 63.625 191.515 63.915 191.560 ;
        RECT 66.000 191.515 66.140 191.670 ;
        RECT 63.625 191.375 66.140 191.515 ;
        RECT 68.760 191.515 68.900 192.055 ;
        RECT 71.445 192.055 73.960 192.195 ;
        RECT 71.445 192.010 71.735 192.055 ;
        RECT 69.130 191.855 69.450 191.915 ;
        RECT 69.605 191.855 69.895 191.900 ;
        RECT 69.130 191.715 69.895 191.855 ;
        RECT 69.130 191.655 69.450 191.715 ;
        RECT 69.605 191.670 69.895 191.715 ;
        RECT 70.510 191.855 70.830 191.915 ;
        RECT 70.985 191.855 71.275 191.900 ;
        RECT 70.510 191.715 71.275 191.855 ;
        RECT 70.510 191.655 70.830 191.715 ;
        RECT 70.985 191.670 71.275 191.715 ;
        RECT 71.890 191.655 72.210 191.915 ;
        RECT 73.820 191.900 73.960 192.055 ;
        RECT 76.505 192.010 76.795 192.240 ;
        RECT 77.040 192.195 77.180 192.335 ;
        RECT 77.425 192.195 77.715 192.240 ;
        RECT 79.250 192.195 79.570 192.255 ;
        RECT 82.100 192.195 82.240 192.395 ;
        RECT 83.850 192.335 84.170 192.395 ;
        RECT 89.000 192.395 97.970 192.535 ;
        RECT 77.040 192.055 77.715 192.195 ;
        RECT 77.425 192.010 77.715 192.055 ;
        RECT 77.960 192.055 79.570 192.195 ;
        RECT 72.365 191.670 72.655 191.900 ;
        RECT 73.745 191.670 74.035 191.900 ;
        RECT 76.965 191.855 77.255 191.900 ;
        RECT 77.960 191.855 78.100 192.055 ;
        RECT 79.250 191.995 79.570 192.055 ;
        RECT 79.800 192.055 82.240 192.195 ;
        RECT 76.965 191.715 78.100 191.855 ;
        RECT 78.790 191.855 79.110 191.915 ;
        RECT 79.800 191.855 79.940 192.055 ;
        RECT 78.790 191.715 79.940 191.855 ;
        RECT 76.965 191.670 77.255 191.715 ;
        RECT 71.980 191.515 72.120 191.655 ;
        RECT 68.760 191.375 72.120 191.515 ;
        RECT 72.440 191.515 72.580 191.670 ;
        RECT 78.790 191.655 79.110 191.715 ;
        RECT 80.170 191.655 80.490 191.915 ;
        RECT 82.100 191.900 82.240 192.055 ;
        RECT 82.485 192.195 82.775 192.240 ;
        RECT 82.485 192.055 83.620 192.195 ;
        RECT 82.485 192.010 82.775 192.055 ;
        RECT 80.645 191.670 80.935 191.900 ;
        RECT 82.025 191.670 82.315 191.900 ;
        RECT 78.330 191.515 78.650 191.575 ;
        RECT 72.440 191.375 78.650 191.515 ;
        RECT 63.625 191.330 63.915 191.375 ;
        RECT 78.330 191.315 78.650 191.375 ;
        RECT 79.710 191.315 80.030 191.575 ;
        RECT 80.720 191.515 80.860 191.670 ;
        RECT 82.930 191.655 83.250 191.915 ;
        RECT 83.480 191.900 83.620 192.055 ;
        RECT 83.405 191.670 83.695 191.900 ;
        RECT 87.070 191.655 87.390 191.915 ;
        RECT 87.545 191.855 87.835 191.900 ;
        RECT 87.990 191.855 88.310 191.915 ;
        RECT 89.000 191.900 89.140 192.395 ;
        RECT 94.430 192.335 94.750 192.395 ;
        RECT 97.650 192.335 97.970 192.395 ;
        RECT 102.800 192.395 105.010 192.535 ;
        RECT 108.805 192.535 109.095 192.580 ;
        RECT 111.925 192.535 112.215 192.580 ;
        RECT 113.815 192.535 114.105 192.580 ;
        RECT 116.510 192.535 116.830 192.595 ;
        RECT 108.805 192.395 114.105 192.535 ;
        RECT 95.810 191.995 96.130 192.255 ;
        RECT 96.285 192.195 96.575 192.240 ;
        RECT 102.250 192.195 102.570 192.255 ;
        RECT 96.285 192.055 102.570 192.195 ;
        RECT 96.285 192.010 96.575 192.055 ;
        RECT 102.250 191.995 102.570 192.055 ;
        RECT 87.545 191.715 88.310 191.855 ;
        RECT 87.545 191.670 87.835 191.715 ;
        RECT 87.990 191.655 88.310 191.715 ;
        RECT 88.925 191.670 89.215 191.900 ;
        RECT 89.370 191.655 89.690 191.915 ;
        RECT 92.590 191.655 92.910 191.915 ;
        RECT 95.365 191.670 95.655 191.900 ;
        RECT 80.720 191.375 85.000 191.515 ;
        RECT 47.510 191.175 47.830 191.235 ;
        RECT 46.680 191.035 47.830 191.175 ;
        RECT 31.410 190.975 31.730 191.035 ;
        RECT 45.225 190.990 45.515 191.035 ;
        RECT 46.130 190.975 46.450 191.035 ;
        RECT 47.510 190.975 47.830 191.035 ;
        RECT 51.650 190.975 51.970 191.235 ;
        RECT 54.410 190.975 54.730 191.235 ;
        RECT 55.330 191.175 55.650 191.235 ;
        RECT 59.485 191.175 59.775 191.220 ;
        RECT 55.330 191.035 59.775 191.175 ;
        RECT 55.330 190.975 55.650 191.035 ;
        RECT 59.485 190.990 59.775 191.035 ;
        RECT 60.390 190.975 60.710 191.235 ;
        RECT 62.230 190.975 62.550 191.235 ;
        RECT 64.530 191.175 64.850 191.235 ;
        RECT 66.845 191.175 67.135 191.220 ;
        RECT 64.530 191.035 67.135 191.175 ;
        RECT 64.530 190.975 64.850 191.035 ;
        RECT 66.845 190.990 67.135 191.035 ;
        RECT 73.730 191.175 74.050 191.235 ;
        RECT 74.665 191.175 74.955 191.220 ;
        RECT 73.730 191.035 74.955 191.175 ;
        RECT 73.730 190.975 74.050 191.035 ;
        RECT 74.665 190.990 74.955 191.035 ;
        RECT 82.930 191.175 83.250 191.235 ;
        RECT 84.325 191.175 84.615 191.220 ;
        RECT 82.930 191.035 84.615 191.175 ;
        RECT 84.860 191.175 85.000 191.375 ;
        RECT 88.450 191.315 88.770 191.575 ;
        RECT 89.830 191.515 90.150 191.575 ;
        RECT 95.440 191.515 95.580 191.670 ;
        RECT 97.650 191.655 97.970 191.915 ;
        RECT 99.490 191.655 99.810 191.915 ;
        RECT 102.800 191.855 102.940 192.395 ;
        RECT 108.805 192.350 109.095 192.395 ;
        RECT 111.925 192.350 112.215 192.395 ;
        RECT 113.815 192.350 114.105 192.395 ;
        RECT 114.760 192.395 116.830 192.535 ;
        RECT 104.550 191.995 104.870 192.255 ;
        RECT 114.760 192.240 114.900 192.395 ;
        RECT 116.510 192.335 116.830 192.395 ;
        RECT 119.820 192.395 124.560 192.535 ;
        RECT 114.685 192.010 114.975 192.240 ;
        RECT 119.270 192.195 119.590 192.255 ;
        RECT 116.600 192.055 119.590 192.195 ;
        RECT 100.040 191.715 102.940 191.855 ;
        RECT 89.830 191.375 95.580 191.515 ;
        RECT 89.830 191.315 90.150 191.375 ;
        RECT 98.585 191.330 98.875 191.560 ;
        RECT 89.370 191.175 89.690 191.235 ;
        RECT 84.860 191.035 89.690 191.175 ;
        RECT 82.930 190.975 83.250 191.035 ;
        RECT 84.325 190.990 84.615 191.035 ;
        RECT 89.370 190.975 89.690 191.035 ;
        RECT 92.130 191.175 92.450 191.235 ;
        RECT 93.525 191.175 93.815 191.220 ;
        RECT 92.130 191.035 93.815 191.175 ;
        RECT 92.130 190.975 92.450 191.035 ;
        RECT 93.525 190.990 93.815 191.035 ;
        RECT 93.970 191.175 94.290 191.235 ;
        RECT 98.660 191.175 98.800 191.330 ;
        RECT 99.030 191.315 99.350 191.575 ;
        RECT 100.040 191.175 100.180 191.715 ;
        RECT 103.170 191.655 103.490 191.915 ;
        RECT 105.010 191.855 105.330 191.915 ;
        RECT 116.600 191.900 116.740 192.055 ;
        RECT 119.270 191.995 119.590 192.055 ;
        RECT 107.725 191.855 108.015 191.875 ;
        RECT 105.010 191.715 108.015 191.855 ;
        RECT 105.010 191.655 105.330 191.715 ;
        RECT 107.725 191.560 108.015 191.715 ;
        RECT 108.805 191.855 109.095 191.900 ;
        RECT 112.385 191.855 112.675 191.900 ;
        RECT 114.220 191.855 114.510 191.900 ;
        RECT 108.805 191.715 114.510 191.855 ;
        RECT 108.805 191.670 109.095 191.715 ;
        RECT 112.385 191.670 112.675 191.715 ;
        RECT 114.220 191.670 114.510 191.715 ;
        RECT 116.525 191.670 116.815 191.900 ;
        RECT 117.445 191.670 117.735 191.900 ;
        RECT 119.820 191.855 119.960 192.395 ;
        RECT 120.190 192.195 120.510 192.255 ;
        RECT 123.425 192.195 123.715 192.240 ;
        RECT 120.190 192.055 123.715 192.195 ;
        RECT 124.420 192.195 124.560 192.395 ;
        RECT 125.250 192.335 125.570 192.595 ;
        RECT 125.710 192.535 126.030 192.595 ;
        RECT 131.230 192.535 131.550 192.595 ;
        RECT 125.710 192.395 131.550 192.535 ;
        RECT 125.710 192.335 126.030 192.395 ;
        RECT 131.230 192.335 131.550 192.395 ;
        RECT 132.610 192.535 132.930 192.595 ;
        RECT 137.670 192.535 137.990 192.595 ;
        RECT 132.610 192.395 137.990 192.535 ;
        RECT 132.610 192.335 132.930 192.395 ;
        RECT 128.930 192.195 129.250 192.255 ;
        RECT 124.420 192.055 129.250 192.195 ;
        RECT 120.190 191.995 120.510 192.055 ;
        RECT 121.660 191.900 121.800 192.055 ;
        RECT 123.425 192.010 123.715 192.055 ;
        RECT 128.930 191.995 129.250 192.055 ;
        RECT 133.990 192.195 134.310 192.255 ;
        RECT 136.305 192.195 136.595 192.240 ;
        RECT 133.990 192.055 136.595 192.195 ;
        RECT 133.990 191.995 134.310 192.055 ;
        RECT 136.305 192.010 136.595 192.055 ;
        RECT 137.300 192.195 137.440 192.395 ;
        RECT 137.670 192.335 137.990 192.395 ;
        RECT 139.065 192.195 139.355 192.240 ;
        RECT 137.300 192.055 139.355 192.195 ;
        RECT 120.665 191.855 120.955 191.900 ;
        RECT 119.820 191.715 120.955 191.855 ;
        RECT 120.665 191.670 120.955 191.715 ;
        RECT 121.585 191.670 121.875 191.900 ;
        RECT 107.425 191.515 108.015 191.560 ;
        RECT 110.665 191.515 111.315 191.560 ;
        RECT 100.500 191.375 106.620 191.515 ;
        RECT 100.500 191.220 100.640 191.375 ;
        RECT 93.970 191.035 100.180 191.175 ;
        RECT 93.970 190.975 94.290 191.035 ;
        RECT 100.425 190.990 100.715 191.220 ;
        RECT 101.330 191.175 101.650 191.235 ;
        RECT 102.265 191.175 102.555 191.220 ;
        RECT 101.330 191.035 102.555 191.175 ;
        RECT 106.480 191.175 106.620 191.375 ;
        RECT 107.425 191.375 111.315 191.515 ;
        RECT 107.425 191.330 107.715 191.375 ;
        RECT 110.665 191.330 111.315 191.375 ;
        RECT 113.305 191.330 113.595 191.560 ;
        RECT 115.130 191.515 115.450 191.575 ;
        RECT 117.520 191.515 117.660 191.670 ;
        RECT 122.950 191.655 123.270 191.915 ;
        RECT 127.565 191.670 127.855 191.900 ;
        RECT 115.130 191.375 117.660 191.515 ;
        RECT 113.380 191.175 113.520 191.330 ;
        RECT 115.130 191.315 115.450 191.375 ;
        RECT 121.110 191.315 121.430 191.575 ;
        RECT 122.275 191.330 122.565 191.560 ;
        RECT 127.640 191.515 127.780 191.670 ;
        RECT 128.010 191.655 128.330 191.915 ;
        RECT 128.470 191.855 128.790 191.915 ;
        RECT 130.325 191.855 130.615 191.900 ;
        RECT 128.470 191.715 130.615 191.855 ;
        RECT 128.470 191.655 128.790 191.715 ;
        RECT 130.325 191.670 130.615 191.715 ;
        RECT 134.450 191.655 134.770 191.915 ;
        RECT 134.925 191.855 135.215 191.900 ;
        RECT 135.370 191.855 135.690 191.915 ;
        RECT 134.925 191.715 135.690 191.855 ;
        RECT 134.925 191.670 135.215 191.715 ;
        RECT 135.370 191.655 135.690 191.715 ;
        RECT 135.830 191.655 136.150 191.915 ;
        RECT 137.300 191.900 137.440 192.055 ;
        RECT 139.065 192.010 139.355 192.055 ;
        RECT 139.600 192.055 141.580 192.195 ;
        RECT 137.225 191.670 137.515 191.900 ;
        RECT 139.600 191.855 139.740 192.055 ;
        RECT 137.760 191.715 139.740 191.855 ;
        RECT 139.985 191.855 140.275 191.900 ;
        RECT 140.890 191.855 141.210 191.915 ;
        RECT 141.440 191.900 141.580 192.055 ;
        RECT 139.985 191.715 141.210 191.855 ;
        RECT 135.920 191.515 136.060 191.655 ;
        RECT 137.760 191.515 137.900 191.715 ;
        RECT 139.985 191.670 140.275 191.715 ;
        RECT 140.890 191.655 141.210 191.715 ;
        RECT 141.365 191.670 141.655 191.900 ;
        RECT 142.270 191.655 142.590 191.915 ;
        RECT 127.640 191.375 135.600 191.515 ;
        RECT 135.920 191.375 137.900 191.515 ;
        RECT 138.145 191.515 138.435 191.560 ;
        RECT 144.125 191.515 144.415 191.560 ;
        RECT 138.145 191.375 144.415 191.515 ;
        RECT 106.480 191.035 113.520 191.175 ;
        RECT 113.750 191.175 114.070 191.235 ;
        RECT 119.745 191.175 120.035 191.220 ;
        RECT 113.750 191.035 120.035 191.175 ;
        RECT 122.350 191.175 122.490 191.330 ;
        RECT 125.710 191.175 126.030 191.235 ;
        RECT 122.350 191.035 126.030 191.175 ;
        RECT 101.330 190.975 101.650 191.035 ;
        RECT 102.265 190.990 102.555 191.035 ;
        RECT 113.750 190.975 114.070 191.035 ;
        RECT 119.745 190.990 120.035 191.035 ;
        RECT 125.710 190.975 126.030 191.035 ;
        RECT 129.390 191.175 129.710 191.235 ;
        RECT 131.245 191.175 131.535 191.220 ;
        RECT 129.390 191.035 131.535 191.175 ;
        RECT 129.390 190.975 129.710 191.035 ;
        RECT 131.245 190.990 131.535 191.035 ;
        RECT 133.070 191.175 133.390 191.235 ;
        RECT 135.460 191.220 135.600 191.375 ;
        RECT 138.145 191.330 138.435 191.375 ;
        RECT 144.125 191.330 144.415 191.375 ;
        RECT 145.965 191.515 146.255 191.560 ;
        RECT 147.330 191.515 147.650 191.575 ;
        RECT 145.965 191.375 147.650 191.515 ;
        RECT 145.965 191.330 146.255 191.375 ;
        RECT 147.330 191.315 147.650 191.375 ;
        RECT 133.545 191.175 133.835 191.220 ;
        RECT 133.070 191.035 133.835 191.175 ;
        RECT 133.070 190.975 133.390 191.035 ;
        RECT 133.545 190.990 133.835 191.035 ;
        RECT 135.385 190.990 135.675 191.220 ;
        RECT 141.810 190.975 142.130 191.235 ;
        RECT 13.860 190.355 147.720 190.835 ;
        RECT 19.910 190.155 20.230 190.215 ;
        RECT 38.770 190.155 39.090 190.215 ;
        RECT 62.230 190.155 62.550 190.215 ;
        RECT 19.910 190.015 34.860 190.155 ;
        RECT 19.910 189.955 20.230 190.015 ;
        RECT 16.690 189.815 17.010 189.875 ;
        RECT 34.720 189.815 34.860 190.015 ;
        RECT 38.770 190.015 62.550 190.155 ;
        RECT 38.770 189.955 39.090 190.015 ;
        RECT 62.230 189.955 62.550 190.015 ;
        RECT 66.830 190.155 67.150 190.215 ;
        RECT 79.710 190.155 80.030 190.215 ;
        RECT 88.450 190.155 88.770 190.215 ;
        RECT 93.970 190.155 94.290 190.215 ;
        RECT 66.830 190.015 94.290 190.155 ;
        RECT 66.830 189.955 67.150 190.015 ;
        RECT 79.710 189.955 80.030 190.015 ;
        RECT 88.450 189.955 88.770 190.015 ;
        RECT 93.970 189.955 94.290 190.015 ;
        RECT 103.630 190.155 103.950 190.215 ;
        RECT 125.250 190.155 125.570 190.215 ;
        RECT 143.650 190.155 143.970 190.215 ;
        RECT 103.630 190.015 118.810 190.155 ;
        RECT 103.630 189.955 103.950 190.015 ;
        RECT 47.050 189.815 47.370 189.875 ;
        RECT 16.690 189.675 22.210 189.815 ;
        RECT 34.720 189.675 47.370 189.815 ;
        RECT 16.690 189.615 17.010 189.675 ;
        RECT 22.070 189.475 22.210 189.675 ;
        RECT 47.050 189.615 47.370 189.675 ;
        RECT 47.510 189.815 47.830 189.875 ;
        RECT 71.430 189.815 71.750 189.875 ;
        RECT 47.510 189.675 71.750 189.815 ;
        RECT 47.510 189.615 47.830 189.675 ;
        RECT 71.430 189.615 71.750 189.675 ;
        RECT 36.470 189.475 36.790 189.535 ;
        RECT 113.750 189.475 114.070 189.535 ;
        RECT 22.070 189.335 34.860 189.475 ;
        RECT 20.370 189.135 20.690 189.195 ;
        RECT 34.720 189.135 34.860 189.335 ;
        RECT 36.470 189.335 114.070 189.475 ;
        RECT 118.670 189.475 118.810 190.015 ;
        RECT 125.250 190.015 143.970 190.155 ;
        RECT 125.250 189.955 125.570 190.015 ;
        RECT 143.650 189.955 143.970 190.015 ;
        RECT 119.270 189.815 119.590 189.875 ;
        RECT 141.810 189.815 142.130 189.875 ;
        RECT 119.270 189.675 142.130 189.815 ;
        RECT 119.270 189.615 119.590 189.675 ;
        RECT 141.810 189.615 142.130 189.675 ;
        RECT 135.830 189.475 136.150 189.535 ;
        RECT 118.670 189.335 136.150 189.475 ;
        RECT 36.470 189.275 36.790 189.335 ;
        RECT 113.750 189.275 114.070 189.335 ;
        RECT 135.830 189.275 136.150 189.335 ;
        RECT 61.770 189.135 62.090 189.195 ;
        RECT 20.370 188.995 33.940 189.135 ;
        RECT 34.720 188.995 62.090 189.135 ;
        RECT 20.370 188.935 20.690 188.995 ;
        RECT 19.450 188.785 19.770 188.845 ;
        RECT 19.450 188.645 31.860 188.785 ;
        RECT 19.450 188.585 19.770 188.645 ;
        RECT 31.720 187.735 31.860 188.645 ;
        RECT 33.800 188.455 33.940 188.995 ;
        RECT 61.770 188.935 62.090 188.995 ;
        RECT 89.370 189.135 89.690 189.195 ;
        RECT 99.490 189.135 99.810 189.195 ;
        RECT 121.110 189.135 121.430 189.195 ;
        RECT 89.370 188.995 121.430 189.135 ;
        RECT 89.370 188.935 89.690 188.995 ;
        RECT 99.490 188.935 99.810 188.995 ;
        RECT 121.110 188.935 121.430 188.995 ;
        RECT 53.950 188.795 54.270 188.855 ;
        RECT 144.110 188.795 144.430 188.855 ;
        RECT 53.950 188.655 144.430 188.795 ;
        RECT 53.950 188.595 54.270 188.655 ;
        RECT 144.110 188.595 144.430 188.655 ;
        RECT 51.190 188.455 51.510 188.515 ;
        RECT 33.800 188.315 51.510 188.455 ;
        RECT 51.190 188.255 51.510 188.315 ;
        RECT 58.090 188.455 58.410 188.515 ;
        RECT 139.510 188.455 139.830 188.465 ;
        RECT 58.090 188.315 139.830 188.455 ;
        RECT 58.090 188.255 58.410 188.315 ;
        RECT 139.510 188.205 139.830 188.315 ;
        RECT 32.330 188.095 32.650 188.155 ;
        RECT 34.630 188.095 34.950 188.155 ;
        RECT 32.330 187.955 34.950 188.095 ;
        RECT 32.330 187.895 32.650 187.955 ;
        RECT 34.630 187.895 34.950 187.955 ;
        RECT 55.790 188.115 56.110 188.175 ;
        RECT 60.390 188.115 60.710 188.175 ;
        RECT 55.790 187.975 60.710 188.115 ;
        RECT 55.790 187.915 56.110 187.975 ;
        RECT 60.390 187.915 60.710 187.975 ;
        RECT 118.810 188.065 119.130 188.125 ;
        RECT 142.270 188.065 142.590 188.125 ;
        RECT 118.810 187.925 142.590 188.065 ;
        RECT 118.810 187.865 119.130 187.925 ;
        RECT 142.270 187.865 142.590 187.925 ;
        RECT 93.510 187.735 93.830 187.795 ;
        RECT 31.720 187.595 93.830 187.735 ;
        RECT 110.490 187.665 110.890 187.790 ;
        RECT 23.090 187.415 23.490 187.540 ;
        RECT 93.510 187.535 93.830 187.595 ;
        RECT 107.040 187.515 110.890 187.665 ;
        RECT 23.090 187.265 27.040 187.415 ;
        RECT 23.090 187.240 23.490 187.265 ;
        RECT 13.890 186.940 14.290 187.240 ;
        RECT 18.490 187.065 18.890 187.240 ;
        RECT 18.490 186.940 26.730 187.065 ;
        RECT 14.040 186.765 14.190 186.940 ;
        RECT 18.615 186.915 26.730 186.940 ;
        RECT 14.040 186.615 26.365 186.765 ;
        RECT 10.365 186.315 26.065 186.465 ;
        RECT 9.915 185.990 25.690 186.140 ;
        RECT 9.615 185.690 25.315 185.840 ;
        RECT 9.315 185.390 24.940 185.540 ;
        RECT 9.015 185.090 24.560 185.240 ;
        RECT 8.715 184.790 24.190 184.940 ;
        RECT 8.415 184.490 23.815 184.640 ;
        RECT 8.115 184.190 23.440 184.340 ;
        RECT 7.815 183.890 23.060 184.040 ;
        RECT 7.515 183.590 22.690 183.740 ;
        RECT 7.215 183.290 22.315 183.440 ;
        RECT 6.915 182.990 21.940 183.140 ;
        RECT 6.615 182.565 7.515 182.715 ;
        RECT 6.315 182.265 7.140 182.415 ;
        RECT 6.015 181.965 6.765 182.115 ;
        RECT 5.715 181.665 6.390 181.810 ;
        RECT 5.415 181.365 6.015 181.515 ;
        RECT 5.115 181.065 5.640 181.215 ;
        RECT 4.815 180.765 5.265 180.915 ;
        RECT 4.515 180.465 4.890 180.615 ;
        RECT 4.215 180.165 4.515 180.315 ;
        RECT 3.915 179.815 4.140 180.015 ;
        RECT 3.990 168.680 4.140 179.815 ;
        RECT 4.365 170.355 4.515 180.165 ;
        RECT 4.740 171.510 4.890 180.465 ;
        RECT 5.115 173.515 5.265 180.765 ;
        RECT 5.490 174.120 5.640 181.065 ;
        RECT 5.865 175.795 6.015 181.365 ;
        RECT 6.245 176.645 6.390 181.665 ;
        RECT 6.615 178.955 6.765 181.965 ;
        RECT 6.990 179.755 7.140 182.265 ;
        RECT 7.365 182.085 7.515 182.565 ;
        RECT 8.035 182.335 21.375 182.815 ;
        RECT 7.290 181.685 7.590 182.085 ;
        RECT 8.790 182.045 21.215 182.195 ;
        RECT 8.155 181.595 8.525 181.625 ;
        RECT 8.065 181.315 8.525 181.595 ;
        RECT 8.790 181.575 8.940 182.045 ;
        RECT 18.215 181.795 18.530 181.860 ;
        RECT 8.065 181.295 8.465 181.315 ;
        RECT 8.705 181.265 9.075 181.575 ;
        RECT 18.215 181.495 18.615 181.795 ;
        RECT 18.215 181.440 18.530 181.495 ;
        RECT 19.005 181.265 19.375 181.575 ;
        RECT 10.855 180.895 11.225 181.125 ;
        RECT 7.290 180.485 7.590 180.885 ;
        RECT 6.915 179.355 7.215 179.755 ;
        RECT 6.540 178.555 6.840 178.955 ;
        RECT 6.915 177.905 7.215 178.305 ;
        RECT 6.540 177.305 6.840 177.705 ;
        RECT 6.170 176.245 6.470 176.645 ;
        RECT 5.790 175.395 6.090 175.795 ;
        RECT 6.170 174.880 6.470 175.280 ;
        RECT 5.790 174.360 6.090 174.760 ;
        RECT 5.420 173.720 5.720 174.120 ;
        RECT 5.040 173.115 5.340 173.515 ;
        RECT 5.420 172.465 5.720 172.865 ;
        RECT 5.040 171.865 5.340 172.265 ;
        RECT 4.745 171.205 4.890 171.510 ;
        RECT 4.670 170.805 4.970 171.205 ;
        RECT 4.290 169.955 4.590 170.355 ;
        RECT 4.670 169.440 4.970 169.840 ;
        RECT 4.290 168.920 4.590 169.320 ;
        RECT 3.920 168.280 4.220 168.680 ;
        RECT 3.540 167.675 3.840 168.075 ;
        RECT 3.920 167.025 4.220 167.425 ;
        RECT 3.540 166.425 3.840 166.825 ;
        RECT 3.615 143.565 3.765 166.425 ;
        RECT 3.990 166.065 4.140 167.025 ;
        RECT 3.915 165.815 4.140 166.065 ;
        RECT 3.915 144.015 4.065 165.815 ;
        RECT 4.365 165.665 4.515 168.920 ;
        RECT 4.215 165.515 4.515 165.665 ;
        RECT 4.215 144.465 4.365 165.515 ;
        RECT 4.740 165.365 4.890 169.440 ;
        RECT 4.515 165.215 4.890 165.365 ;
        RECT 4.515 144.915 4.665 165.215 ;
        RECT 5.115 165.065 5.265 171.865 ;
        RECT 4.815 164.915 5.265 165.065 ;
        RECT 4.815 145.365 4.965 164.915 ;
        RECT 5.490 164.765 5.640 172.465 ;
        RECT 5.115 164.615 5.640 164.765 ;
        RECT 5.115 145.815 5.265 164.615 ;
        RECT 5.865 164.465 6.015 174.360 ;
        RECT 5.415 164.315 6.015 164.465 ;
        RECT 5.415 146.265 5.565 164.315 ;
        RECT 6.245 164.165 6.390 174.880 ;
        RECT 5.715 164.020 6.390 164.165 ;
        RECT 5.715 164.015 6.365 164.020 ;
        RECT 5.715 147.165 5.865 164.015 ;
        RECT 6.615 163.865 6.765 177.305 ;
        RECT 6.015 163.715 6.765 163.865 ;
        RECT 6.015 147.615 6.165 163.715 ;
        RECT 6.990 163.565 7.140 177.905 ;
        RECT 6.315 163.415 7.140 163.565 ;
        RECT 6.315 148.065 6.465 163.415 ;
        RECT 7.365 163.265 7.515 180.485 ;
        RECT 10.815 180.395 11.265 180.895 ;
        RECT 19.090 180.395 19.240 181.265 ;
        RECT 21.065 181.245 21.215 182.045 ;
        RECT 20.915 181.225 21.315 181.245 ;
        RECT 20.905 180.945 21.315 181.225 ;
        RECT 20.905 180.915 21.275 180.945 ;
        RECT 10.815 180.245 19.240 180.395 ;
        RECT 8.035 179.615 21.375 180.095 ;
        RECT 8.115 179.145 8.515 179.445 ;
        RECT 10.940 179.315 19.240 179.465 ;
        RECT 8.215 178.725 8.365 179.145 ;
        RECT 10.940 178.925 11.090 179.315 ;
        RECT 8.105 178.415 8.475 178.725 ;
        RECT 10.855 178.615 11.225 178.925 ;
        RECT 14.055 178.865 14.425 178.895 ;
        RECT 14.015 178.815 14.425 178.865 ;
        RECT 18.215 178.845 18.615 179.145 ;
        RECT 14.015 178.665 16.065 178.815 ;
        RECT 8.705 178.135 9.075 178.445 ;
        RECT 10.915 178.245 11.065 178.615 ;
        RECT 14.015 178.585 14.425 178.665 ;
        RECT 14.015 178.565 14.415 178.585 ;
        RECT 11.315 178.445 11.715 178.465 ;
        RECT 15.915 178.445 16.065 178.665 ;
        RECT 8.790 177.665 8.940 178.135 ;
        RECT 10.765 177.945 11.165 178.245 ;
        RECT 11.315 178.165 11.725 178.445 ;
        RECT 11.355 178.135 11.725 178.165 ;
        RECT 11.905 178.135 12.275 178.445 ;
        RECT 14.955 178.415 15.325 178.445 ;
        RECT 14.955 178.135 15.365 178.415 ;
        RECT 15.805 178.135 16.175 178.445 ;
        RECT 17.675 178.195 18.045 178.445 ;
        RECT 17.615 178.135 18.045 178.195 ;
        RECT 18.315 178.180 18.465 178.845 ;
        RECT 19.090 178.445 19.240 179.315 ;
        RECT 20.905 178.465 21.275 178.495 ;
        RECT 12.015 177.955 12.165 178.135 ;
        RECT 14.965 178.115 15.365 178.135 ;
        RECT 17.615 177.955 18.015 178.135 ;
        RECT 12.015 177.895 18.015 177.955 ;
        RECT 12.015 177.805 17.910 177.895 ;
        RECT 18.185 177.870 18.555 178.180 ;
        RECT 19.005 178.135 19.375 178.445 ;
        RECT 20.905 178.185 21.315 178.465 ;
        RECT 20.915 178.165 21.315 178.185 ;
        RECT 21.065 177.665 21.215 178.165 ;
        RECT 8.790 177.515 21.215 177.665 ;
        RECT 8.035 176.895 21.375 177.375 ;
        RECT 8.790 176.605 21.215 176.755 ;
        RECT 8.155 176.155 8.525 176.185 ;
        RECT 8.065 175.875 8.525 176.155 ;
        RECT 8.790 176.135 8.940 176.605 ;
        RECT 12.015 176.315 17.940 176.465 ;
        RECT 12.015 176.135 12.165 176.315 ;
        RECT 14.965 176.135 15.365 176.155 ;
        RECT 17.790 176.135 17.940 176.315 ;
        RECT 18.215 176.355 18.530 176.420 ;
        RECT 8.065 175.855 8.465 175.875 ;
        RECT 8.705 175.825 9.075 176.135 ;
        RECT 11.355 176.105 11.725 176.135 ;
        RECT 11.315 175.825 11.725 176.105 ;
        RECT 11.905 175.825 12.275 176.135 ;
        RECT 14.955 175.855 15.365 176.135 ;
        RECT 14.955 175.825 15.325 175.855 ;
        RECT 15.805 175.825 16.175 176.135 ;
        RECT 17.705 175.825 18.075 176.135 ;
        RECT 18.215 176.055 18.615 176.355 ;
        RECT 18.215 176.000 18.530 176.055 ;
        RECT 19.005 175.825 19.375 176.135 ;
        RECT 11.315 175.805 11.715 175.825 ;
        RECT 14.015 175.685 14.415 175.705 ;
        RECT 10.855 175.455 11.225 175.685 ;
        RECT 14.015 175.605 14.425 175.685 ;
        RECT 15.915 175.605 16.065 175.825 ;
        RECT 14.015 175.455 16.065 175.605 ;
        RECT 10.815 174.955 11.265 175.455 ;
        RECT 14.015 175.405 14.425 175.455 ;
        RECT 17.790 175.405 17.940 175.825 ;
        RECT 14.055 175.375 14.425 175.405 ;
        RECT 17.665 175.105 18.065 175.405 ;
        RECT 19.090 174.955 19.240 175.825 ;
        RECT 21.065 175.805 21.215 176.605 ;
        RECT 20.915 175.785 21.315 175.805 ;
        RECT 20.905 175.505 21.315 175.785 ;
        RECT 20.905 175.475 21.275 175.505 ;
        RECT 10.815 174.805 19.240 174.955 ;
        RECT 8.035 174.175 21.375 174.655 ;
        RECT 8.115 173.705 8.515 174.005 ;
        RECT 10.940 173.875 19.240 174.025 ;
        RECT 8.215 173.285 8.365 173.705 ;
        RECT 10.940 173.485 11.090 173.875 ;
        RECT 8.105 172.975 8.475 173.285 ;
        RECT 10.855 173.175 11.225 173.485 ;
        RECT 14.055 173.425 14.425 173.455 ;
        RECT 14.015 173.375 14.425 173.425 ;
        RECT 18.215 173.405 18.615 173.705 ;
        RECT 14.015 173.225 16.065 173.375 ;
        RECT 8.705 172.695 9.075 173.005 ;
        RECT 10.915 172.805 11.065 173.175 ;
        RECT 14.015 173.145 14.425 173.225 ;
        RECT 14.015 173.125 14.415 173.145 ;
        RECT 11.315 173.005 11.715 173.025 ;
        RECT 15.915 173.005 16.065 173.225 ;
        RECT 8.790 172.225 8.940 172.695 ;
        RECT 10.765 172.505 11.165 172.805 ;
        RECT 11.315 172.725 11.725 173.005 ;
        RECT 11.355 172.695 11.725 172.725 ;
        RECT 11.905 172.695 12.275 173.005 ;
        RECT 14.955 172.975 15.325 173.005 ;
        RECT 14.955 172.695 15.365 172.975 ;
        RECT 15.805 172.695 16.175 173.005 ;
        RECT 17.675 172.755 18.045 173.005 ;
        RECT 17.615 172.695 18.045 172.755 ;
        RECT 18.315 172.740 18.465 173.405 ;
        RECT 19.090 173.005 19.240 173.875 ;
        RECT 20.905 173.025 21.275 173.055 ;
        RECT 12.015 172.515 12.165 172.695 ;
        RECT 14.965 172.675 15.365 172.695 ;
        RECT 17.615 172.515 18.015 172.695 ;
        RECT 12.015 172.455 18.015 172.515 ;
        RECT 12.015 172.365 17.910 172.455 ;
        RECT 18.185 172.430 18.555 172.740 ;
        RECT 19.005 172.695 19.375 173.005 ;
        RECT 20.905 172.745 21.315 173.025 ;
        RECT 20.915 172.725 21.315 172.745 ;
        RECT 21.065 172.225 21.215 172.725 ;
        RECT 8.790 172.075 21.215 172.225 ;
        RECT 8.035 171.455 21.375 171.935 ;
        RECT 8.790 171.165 21.215 171.315 ;
        RECT 8.155 170.715 8.525 170.745 ;
        RECT 8.065 170.435 8.525 170.715 ;
        RECT 8.790 170.695 8.940 171.165 ;
        RECT 12.015 170.875 17.940 171.025 ;
        RECT 12.015 170.695 12.165 170.875 ;
        RECT 14.965 170.695 15.365 170.715 ;
        RECT 17.790 170.695 17.940 170.875 ;
        RECT 18.215 170.915 18.530 170.980 ;
        RECT 8.065 170.415 8.465 170.435 ;
        RECT 8.705 170.385 9.075 170.695 ;
        RECT 11.355 170.665 11.725 170.695 ;
        RECT 11.315 170.385 11.725 170.665 ;
        RECT 11.905 170.385 12.275 170.695 ;
        RECT 14.955 170.415 15.365 170.695 ;
        RECT 14.955 170.385 15.325 170.415 ;
        RECT 15.805 170.385 16.175 170.695 ;
        RECT 17.705 170.385 18.075 170.695 ;
        RECT 18.215 170.615 18.615 170.915 ;
        RECT 18.215 170.560 18.530 170.615 ;
        RECT 19.005 170.385 19.375 170.695 ;
        RECT 11.315 170.365 11.715 170.385 ;
        RECT 14.015 170.245 14.415 170.265 ;
        RECT 10.855 170.015 11.225 170.245 ;
        RECT 14.015 170.165 14.425 170.245 ;
        RECT 15.915 170.165 16.065 170.385 ;
        RECT 14.015 170.015 16.065 170.165 ;
        RECT 10.815 169.515 11.265 170.015 ;
        RECT 14.015 169.965 14.425 170.015 ;
        RECT 17.790 169.965 17.940 170.385 ;
        RECT 14.055 169.935 14.425 169.965 ;
        RECT 17.665 169.665 18.065 169.965 ;
        RECT 19.090 169.515 19.240 170.385 ;
        RECT 21.065 170.365 21.215 171.165 ;
        RECT 20.915 170.345 21.315 170.365 ;
        RECT 20.905 170.065 21.315 170.345 ;
        RECT 20.905 170.035 21.275 170.065 ;
        RECT 10.815 169.365 19.240 169.515 ;
        RECT 8.035 168.735 21.375 169.215 ;
        RECT 8.115 168.265 8.515 168.565 ;
        RECT 10.940 168.435 19.240 168.585 ;
        RECT 8.215 167.845 8.365 168.265 ;
        RECT 10.940 168.045 11.090 168.435 ;
        RECT 8.105 167.535 8.475 167.845 ;
        RECT 10.855 167.735 11.225 168.045 ;
        RECT 14.055 167.985 14.425 168.015 ;
        RECT 14.015 167.935 14.425 167.985 ;
        RECT 18.215 167.965 18.615 168.265 ;
        RECT 14.015 167.785 16.065 167.935 ;
        RECT 8.705 167.255 9.075 167.565 ;
        RECT 10.915 167.365 11.065 167.735 ;
        RECT 14.015 167.705 14.425 167.785 ;
        RECT 14.015 167.685 14.415 167.705 ;
        RECT 11.315 167.565 11.715 167.585 ;
        RECT 15.915 167.565 16.065 167.785 ;
        RECT 8.790 166.785 8.940 167.255 ;
        RECT 10.765 167.065 11.165 167.365 ;
        RECT 11.315 167.285 11.725 167.565 ;
        RECT 11.355 167.255 11.725 167.285 ;
        RECT 11.905 167.255 12.275 167.565 ;
        RECT 14.955 167.535 15.325 167.565 ;
        RECT 14.955 167.255 15.365 167.535 ;
        RECT 15.805 167.255 16.175 167.565 ;
        RECT 17.675 167.315 18.045 167.565 ;
        RECT 17.615 167.255 18.045 167.315 ;
        RECT 18.315 167.300 18.465 167.965 ;
        RECT 19.090 167.565 19.240 168.435 ;
        RECT 21.790 168.250 21.940 182.990 ;
        RECT 22.165 168.795 22.315 183.290 ;
        RECT 22.540 171.000 22.690 183.590 ;
        RECT 22.915 171.610 23.060 183.890 ;
        RECT 23.290 173.690 23.440 184.190 ;
        RECT 23.665 174.235 23.815 184.490 ;
        RECT 24.040 176.440 24.190 184.790 ;
        RECT 24.415 177.050 24.560 185.090 ;
        RECT 24.790 179.130 24.940 185.390 ;
        RECT 25.165 179.675 25.315 185.690 ;
        RECT 25.540 182.255 25.690 185.990 ;
        RECT 25.465 181.855 25.765 182.255 ;
        RECT 25.465 180.805 25.765 181.205 ;
        RECT 25.090 179.275 25.390 179.675 ;
        RECT 24.715 178.730 25.015 179.130 ;
        RECT 25.090 178.075 25.390 178.475 ;
        RECT 24.715 177.325 25.015 177.725 ;
        RECT 24.415 177.015 24.565 177.050 ;
        RECT 24.340 176.615 24.640 177.015 ;
        RECT 23.965 176.040 24.265 176.440 ;
        RECT 24.340 175.365 24.640 175.765 ;
        RECT 24.415 175.350 24.565 175.365 ;
        RECT 23.965 174.715 24.265 175.115 ;
        RECT 23.590 173.835 23.890 174.235 ;
        RECT 23.215 173.290 23.515 173.690 ;
        RECT 23.590 172.635 23.890 173.035 ;
        RECT 23.215 171.885 23.515 172.285 ;
        RECT 22.915 171.575 23.065 171.610 ;
        RECT 22.840 171.175 23.140 171.575 ;
        RECT 22.465 170.600 22.765 171.000 ;
        RECT 22.840 169.925 23.140 170.325 ;
        RECT 22.915 169.910 23.065 169.925 ;
        RECT 22.465 169.275 22.765 169.675 ;
        RECT 22.090 168.395 22.390 168.795 ;
        RECT 21.715 167.850 22.015 168.250 ;
        RECT 20.905 167.585 21.275 167.615 ;
        RECT 12.015 167.075 12.165 167.255 ;
        RECT 14.965 167.235 15.365 167.255 ;
        RECT 17.615 167.075 18.015 167.255 ;
        RECT 12.015 167.015 18.015 167.075 ;
        RECT 12.015 166.925 17.910 167.015 ;
        RECT 18.185 166.990 18.555 167.300 ;
        RECT 19.005 167.255 19.375 167.565 ;
        RECT 20.905 167.305 21.315 167.585 ;
        RECT 20.915 167.285 21.315 167.305 ;
        RECT 21.065 166.785 21.215 167.285 ;
        RECT 22.090 167.195 22.390 167.595 ;
        RECT 8.790 166.635 21.215 166.785 ;
        RECT 8.035 166.015 21.375 166.495 ;
        RECT 21.715 166.445 22.015 166.845 ;
        RECT 21.790 165.830 21.940 166.445 ;
        RECT 6.615 163.115 7.515 163.265 ;
        RECT 7.665 165.680 21.940 165.830 ;
        RECT 6.615 148.515 6.765 163.115 ;
        RECT 7.665 162.965 7.815 165.680 ;
        RECT 22.165 165.530 22.315 167.195 ;
        RECT 6.915 162.815 7.815 162.965 ;
        RECT 7.965 165.380 22.315 165.530 ;
        RECT 6.915 148.965 7.065 162.815 ;
        RECT 7.965 162.665 8.115 165.380 ;
        RECT 22.540 165.230 22.690 169.275 ;
        RECT 7.215 162.515 8.115 162.665 ;
        RECT 8.265 165.105 22.690 165.230 ;
        RECT 22.915 166.295 23.060 169.910 ;
        RECT 8.265 165.080 22.670 165.105 ;
        RECT 7.215 149.415 7.365 162.515 ;
        RECT 8.265 162.365 8.415 165.080 ;
        RECT 22.915 164.930 23.065 166.295 ;
        RECT 7.515 162.215 8.415 162.365 ;
        RECT 8.565 164.780 23.065 164.930 ;
        RECT 7.515 149.865 7.665 162.215 ;
        RECT 8.565 162.065 8.715 164.780 ;
        RECT 23.290 164.630 23.440 171.885 ;
        RECT 7.815 161.915 8.715 162.065 ;
        RECT 8.865 164.480 23.440 164.630 ;
        RECT 7.815 150.315 7.965 161.915 ;
        RECT 8.865 161.765 9.015 164.480 ;
        RECT 23.665 164.330 23.815 172.635 ;
        RECT 8.115 161.615 9.015 161.765 ;
        RECT 9.165 164.180 23.815 164.330 ;
        RECT 8.115 150.765 8.265 161.615 ;
        RECT 9.165 161.465 9.315 164.180 ;
        RECT 24.040 164.030 24.190 174.715 ;
        RECT 8.415 161.315 9.315 161.465 ;
        RECT 9.465 163.880 24.190 164.030 ;
        RECT 24.415 166.295 24.560 175.350 ;
        RECT 8.415 151.215 8.565 161.315 ;
        RECT 9.465 161.165 9.615 163.880 ;
        RECT 24.415 163.730 24.565 166.295 ;
        RECT 8.715 161.015 9.615 161.165 ;
        RECT 9.765 163.580 24.565 163.730 ;
        RECT 8.715 151.665 8.865 161.015 ;
        RECT 9.765 160.865 9.915 163.580 ;
        RECT 24.790 163.430 24.940 177.325 ;
        RECT 9.015 160.715 9.915 160.865 ;
        RECT 10.065 163.280 24.940 163.430 ;
        RECT 9.015 152.115 9.165 160.715 ;
        RECT 10.065 160.565 10.215 163.280 ;
        RECT 25.165 163.130 25.315 178.075 ;
        RECT 9.315 160.415 10.215 160.565 ;
        RECT 10.365 162.980 25.315 163.130 ;
        RECT 9.315 152.565 9.465 160.415 ;
        RECT 10.365 160.265 10.515 162.980 ;
        RECT 25.540 162.830 25.690 180.805 ;
        RECT 10.670 162.815 25.690 162.830 ;
        RECT 9.615 160.115 10.515 160.265 ;
        RECT 10.665 162.690 25.690 162.815 ;
        RECT 9.615 153.015 9.765 160.115 ;
        RECT 10.665 159.965 10.815 162.690 ;
        RECT 25.915 162.515 26.065 186.315 ;
        RECT 9.915 159.815 10.815 159.965 ;
        RECT 10.965 162.365 26.065 162.515 ;
        RECT 9.915 153.590 10.065 159.815 ;
        RECT 10.965 159.665 11.115 162.365 ;
        RECT 26.215 162.215 26.365 186.615 ;
        RECT 26.580 173.020 26.730 186.915 ;
        RECT 26.890 178.440 27.040 187.265 ;
        RECT 105.890 186.465 106.290 186.640 ;
        RECT 105.890 186.340 106.890 186.465 ;
        RECT 106.015 186.315 106.890 186.340 ;
        RECT 96.640 186.165 97.040 186.240 ;
        RECT 96.640 186.015 106.590 186.165 ;
        RECT 96.640 185.940 97.040 186.015 ;
        RECT 32.290 185.715 32.690 185.790 ;
        RECT 32.290 185.565 106.290 185.715 ;
        RECT 32.290 185.490 32.690 185.565 ;
        RECT 41.440 185.265 41.840 185.340 ;
        RECT 41.440 185.115 105.990 185.265 ;
        RECT 41.440 185.040 41.840 185.115 ;
        RECT 82.890 184.815 83.290 184.890 ;
        RECT 30.765 184.665 83.290 184.815 ;
        RECT 26.890 178.140 27.290 178.440 ;
        RECT 26.505 172.620 26.805 173.020 ;
        RECT 10.365 159.515 11.115 159.665 ;
        RECT 11.265 162.065 30.315 162.215 ;
        RECT 10.365 158.840 10.515 159.515 ;
        RECT 11.265 159.365 11.415 162.065 ;
        RECT 30.165 160.615 30.315 162.065 ;
        RECT 30.765 161.740 30.915 184.665 ;
        RECT 82.890 184.590 83.290 184.665 ;
        RECT 105.240 184.490 105.640 184.790 ;
        RECT 73.690 184.365 74.090 184.440 ;
        RECT 31.065 184.215 74.090 184.365 ;
        RECT 31.065 162.040 31.215 184.215 ;
        RECT 73.690 184.140 74.090 184.215 ;
        RECT 64.490 183.915 64.890 183.990 ;
        RECT 31.365 183.765 64.890 183.915 ;
        RECT 31.365 162.340 31.515 183.765 ;
        RECT 64.490 183.690 64.890 183.765 ;
        RECT 104.790 183.465 105.190 183.540 ;
        RECT 31.665 183.315 105.190 183.465 ;
        RECT 31.665 162.640 31.815 183.315 ;
        RECT 104.790 183.240 105.190 183.315 ;
        RECT 55.240 183.015 55.640 183.040 ;
        RECT 103.340 183.015 103.740 183.090 ;
        RECT 31.965 182.865 55.640 183.015 ;
        RECT 31.965 162.940 32.115 182.865 ;
        RECT 55.240 182.740 55.640 182.865 ;
        RECT 75.465 182.865 103.740 183.015 ;
        RECT 50.690 182.565 51.090 182.590 ;
        RECT 32.265 182.415 51.090 182.565 ;
        RECT 32.265 163.240 32.415 182.415 ;
        RECT 50.690 182.290 51.090 182.415 ;
        RECT 75.465 182.115 75.615 182.865 ;
        RECT 103.340 182.790 103.740 182.865 ;
        RECT 42.565 181.965 75.615 182.115 ;
        RECT 42.565 181.715 42.715 181.965 ;
        RECT 33.290 181.565 42.715 181.715 ;
        RECT 76.090 181.630 78.040 182.690 ;
        RECT 32.565 178.090 32.965 178.390 ;
        RECT 32.590 163.865 32.740 178.090 ;
        RECT 33.290 172.990 33.440 181.565 ;
        RECT 47.420 180.830 71.320 181.630 ;
        RECT 71.870 180.830 102.970 181.630 ;
        RECT 34.640 179.840 46.040 180.640 ;
        RECT 35.590 179.600 39.270 179.840 ;
        RECT 40.180 179.390 40.470 179.410 ;
        RECT 39.440 179.190 40.470 179.390 ;
        RECT 41.760 179.365 42.050 179.410 ;
        RECT 35.580 178.110 36.000 178.470 ;
        RECT 38.590 178.460 38.990 178.490 ;
        RECT 38.570 178.165 39.005 178.460 ;
        RECT 39.440 177.790 39.640 179.190 ;
        RECT 40.180 179.180 40.470 179.190 ;
        RECT 41.040 179.215 42.050 179.365 ;
        RECT 39.990 178.840 40.220 178.975 ;
        RECT 39.840 178.540 40.240 178.840 ;
        RECT 39.990 177.975 40.220 178.540 ;
        RECT 40.430 178.115 40.660 178.975 ;
        RECT 40.430 177.975 40.890 178.115 ;
        RECT 40.515 177.965 40.890 177.975 ;
        RECT 39.390 177.770 40.440 177.790 ;
        RECT 39.390 177.590 40.470 177.770 ;
        RECT 34.640 177.360 36.040 177.440 ;
        RECT 34.640 176.880 39.270 177.360 ;
        RECT 34.640 176.840 36.040 176.880 ;
        RECT 33.190 172.690 33.590 172.990 ;
        RECT 34.640 171.940 35.240 176.840 ;
        RECT 39.440 176.390 39.640 177.590 ;
        RECT 40.180 177.540 40.470 177.590 ;
        RECT 40.740 177.190 40.890 177.965 ;
        RECT 40.490 176.890 40.890 177.190 ;
        RECT 40.180 176.390 40.470 176.410 ;
        RECT 39.390 176.190 40.470 176.390 ;
        RECT 35.580 175.760 36.000 176.120 ;
        RECT 38.590 176.075 38.990 176.090 ;
        RECT 38.560 175.775 39.010 176.075 ;
        RECT 39.440 174.740 39.640 176.190 ;
        RECT 40.180 176.180 40.470 176.190 ;
        RECT 39.990 175.790 40.220 175.975 ;
        RECT 39.840 175.490 40.240 175.790 ;
        RECT 39.990 174.975 40.220 175.490 ;
        RECT 40.430 175.240 40.660 175.975 ;
        RECT 40.430 174.975 40.790 175.240 ;
        RECT 40.180 174.740 40.470 174.770 ;
        RECT 35.590 174.160 39.270 174.640 ;
        RECT 39.440 174.540 40.490 174.740 ;
        RECT 39.440 173.240 39.640 174.540 ;
        RECT 40.640 173.390 40.790 174.975 ;
        RECT 41.040 174.790 41.190 179.215 ;
        RECT 41.760 179.180 42.050 179.215 ;
        RECT 43.340 179.365 43.630 179.410 ;
        RECT 44.920 179.390 45.210 179.410 ;
        RECT 43.340 179.215 44.340 179.365 ;
        RECT 43.340 179.180 43.630 179.215 ;
        RECT 41.570 178.840 41.800 178.975 ;
        RECT 41.440 178.540 41.840 178.840 ;
        RECT 41.570 178.340 41.800 178.540 ;
        RECT 41.440 178.040 41.840 178.340 ;
        RECT 41.570 177.890 41.800 178.040 ;
        RECT 41.440 177.590 41.840 177.890 ;
        RECT 41.570 174.975 41.800 177.590 ;
        RECT 42.010 177.190 42.240 178.975 ;
        RECT 43.150 177.190 43.380 178.975 ;
        RECT 43.590 178.840 43.820 178.975 ;
        RECT 43.540 178.540 43.940 178.840 ;
        RECT 43.590 178.340 43.820 178.540 ;
        RECT 43.540 178.040 43.940 178.340 ;
        RECT 43.590 177.890 43.820 178.040 ;
        RECT 43.540 177.590 43.940 177.890 ;
        RECT 41.940 176.890 42.340 177.190 ;
        RECT 43.040 176.890 43.440 177.190 ;
        RECT 42.010 175.715 42.240 176.890 ;
        RECT 43.150 175.715 43.380 176.890 ;
        RECT 42.010 175.565 42.540 175.715 ;
        RECT 42.010 174.975 42.240 175.565 ;
        RECT 40.940 174.715 41.340 174.790 ;
        RECT 41.760 174.715 42.050 174.770 ;
        RECT 40.940 174.565 42.050 174.715 ;
        RECT 40.940 174.490 41.340 174.565 ;
        RECT 41.760 174.540 42.050 174.565 ;
        RECT 39.440 173.040 40.490 173.240 ;
        RECT 35.645 172.990 36.100 173.025 ;
        RECT 37.190 173.020 37.640 173.040 ;
        RECT 35.640 172.725 36.100 172.990 ;
        RECT 35.640 172.690 36.040 172.725 ;
        RECT 37.180 172.660 37.640 173.020 ;
        RECT 37.190 172.640 37.640 172.660 ;
        RECT 34.640 171.920 36.040 171.940 ;
        RECT 34.640 171.440 38.350 171.920 ;
        RECT 34.640 171.340 36.040 171.440 ;
        RECT 34.640 167.540 35.240 171.340 ;
        RECT 37.240 170.640 37.640 170.740 ;
        RECT 39.470 170.640 39.640 173.040 ;
        RECT 40.185 172.990 40.475 173.040 ;
        RECT 40.640 172.990 40.940 173.390 ;
        RECT 41.140 173.190 41.290 174.490 ;
        RECT 42.390 174.240 42.540 175.565 ;
        RECT 42.840 175.565 43.380 175.715 ;
        RECT 42.840 174.790 42.990 175.565 ;
        RECT 43.150 174.975 43.380 175.565 ;
        RECT 43.590 174.975 43.820 177.590 ;
        RECT 42.740 174.490 43.140 174.790 ;
        RECT 43.340 174.715 43.630 174.770 ;
        RECT 44.190 174.715 44.340 179.215 ;
        RECT 44.890 179.190 45.940 179.390 ;
        RECT 44.920 179.180 45.210 179.190 ;
        RECT 44.730 178.115 44.960 178.975 ;
        RECT 45.170 178.840 45.400 178.975 ;
        RECT 45.140 178.540 45.540 178.840 ;
        RECT 44.490 177.975 44.960 178.115 ;
        RECT 45.170 177.975 45.400 178.540 ;
        RECT 44.490 177.965 44.865 177.975 ;
        RECT 44.490 177.190 44.640 177.965 ;
        RECT 44.920 177.740 45.210 177.770 ;
        RECT 45.740 177.740 45.940 179.190 ;
        RECT 44.890 177.540 45.940 177.740 ;
        RECT 44.490 176.890 44.890 177.190 ;
        RECT 44.920 176.390 45.210 176.410 ;
        RECT 45.740 176.390 45.940 177.540 ;
        RECT 44.890 176.190 45.940 176.390 ;
        RECT 44.920 176.180 45.210 176.190 ;
        RECT 44.730 175.240 44.960 175.975 ;
        RECT 45.170 175.790 45.400 175.975 ;
        RECT 45.140 175.490 45.540 175.790 ;
        RECT 43.340 174.565 44.340 174.715 ;
        RECT 43.340 174.540 43.630 174.565 ;
        RECT 42.240 173.940 42.640 174.240 ;
        RECT 41.765 173.190 42.055 173.220 ;
        RECT 41.140 172.990 42.055 173.190 ;
        RECT 39.995 172.740 40.225 172.830 ;
        RECT 39.890 172.440 40.290 172.740 ;
        RECT 39.995 171.940 40.225 172.440 ;
        RECT 39.890 171.640 40.290 171.940 ;
        RECT 39.995 170.830 40.225 171.640 ;
        RECT 40.435 171.390 40.665 172.830 ;
        RECT 41.140 171.640 41.290 172.990 ;
        RECT 41.575 172.190 41.805 172.830 ;
        RECT 42.015 172.490 42.245 172.830 ;
        RECT 42.390 172.490 42.540 173.940 ;
        RECT 42.015 172.340 42.540 172.490 ;
        RECT 42.840 172.490 42.990 174.490 ;
        RECT 44.190 174.240 44.340 174.565 ;
        RECT 44.590 174.975 44.960 175.240 ;
        RECT 45.170 174.975 45.400 175.490 ;
        RECT 44.040 173.940 44.440 174.240 ;
        RECT 43.345 173.165 43.635 173.220 ;
        RECT 44.090 173.165 44.240 173.940 ;
        RECT 44.590 173.390 44.740 174.975 ;
        RECT 44.920 174.740 45.210 174.770 ;
        RECT 45.740 174.740 45.940 176.190 ;
        RECT 44.890 174.540 45.940 174.740 ;
        RECT 43.345 173.015 44.240 173.165 ;
        RECT 43.345 172.990 43.635 173.015 ;
        RECT 43.155 172.490 43.385 172.830 ;
        RECT 42.840 172.340 43.385 172.490 ;
        RECT 41.440 171.890 41.840 172.190 ;
        RECT 41.575 171.830 41.805 171.890 ;
        RECT 42.015 171.830 42.245 172.340 ;
        RECT 43.155 171.830 43.385 172.340 ;
        RECT 43.595 172.240 43.825 172.830 ;
        RECT 43.595 172.190 43.940 172.240 ;
        RECT 43.590 171.890 43.940 172.190 ;
        RECT 43.595 171.840 43.940 171.890 ;
        RECT 43.595 171.830 43.825 171.840 ;
        RECT 41.765 171.640 42.055 171.670 ;
        RECT 41.140 171.440 42.055 171.640 ;
        RECT 43.345 171.615 43.635 171.670 ;
        RECT 44.090 171.615 44.240 173.015 ;
        RECT 44.440 172.990 44.740 173.390 ;
        RECT 44.925 173.190 45.215 173.220 ;
        RECT 45.740 173.190 45.940 174.540 ;
        RECT 44.925 172.990 45.940 173.190 ;
        RECT 43.345 171.465 44.240 171.615 ;
        RECT 43.345 171.440 43.635 171.465 ;
        RECT 44.090 171.440 44.240 171.465 ;
        RECT 44.735 171.390 44.965 172.830 ;
        RECT 40.435 171.090 40.840 171.390 ;
        RECT 44.490 171.090 44.965 171.390 ;
        RECT 40.435 170.830 40.665 171.090 ;
        RECT 44.735 170.830 44.965 171.090 ;
        RECT 45.175 172.740 45.405 172.830 ;
        RECT 45.175 172.440 45.590 172.740 ;
        RECT 45.175 171.940 45.405 172.440 ;
        RECT 45.175 171.640 45.590 171.940 ;
        RECT 45.175 170.830 45.405 171.640 ;
        RECT 40.185 170.640 40.475 170.670 ;
        RECT 44.925 170.640 45.215 170.670 ;
        RECT 45.790 170.640 45.940 172.990 ;
        RECT 37.240 170.440 45.940 170.640 ;
        RECT 39.890 167.540 40.290 170.240 ;
        RECT 40.440 169.890 40.840 170.190 ;
        RECT 41.440 169.890 41.840 170.190 ;
        RECT 43.590 170.015 43.990 170.190 ;
        RECT 43.540 169.890 43.990 170.015 ;
        RECT 44.490 169.890 44.890 170.190 ;
        RECT 40.640 169.260 40.790 169.890 ;
        RECT 40.940 169.640 41.230 169.650 ;
        RECT 40.940 169.260 41.240 169.640 ;
        RECT 41.640 169.260 41.790 169.890 ;
        RECT 42.990 169.440 43.390 169.740 ;
        RECT 43.040 169.420 43.330 169.440 ;
        RECT 43.540 169.260 43.690 169.890 ;
        RECT 44.490 169.260 44.640 169.890 ;
        RECT 40.640 168.940 41.440 169.260 ;
        RECT 41.640 169.040 42.010 169.260 ;
        RECT 40.730 168.590 40.960 168.940 ;
        RECT 41.210 168.590 41.440 168.940 ;
        RECT 40.730 168.290 41.440 168.590 ;
        RECT 40.730 168.260 40.960 168.290 ;
        RECT 41.210 168.260 41.440 168.290 ;
        RECT 41.780 168.260 42.010 169.040 ;
        RECT 42.260 168.590 42.490 169.260 ;
        RECT 42.830 168.590 43.060 169.260 ;
        RECT 42.260 168.290 43.060 168.590 ;
        RECT 42.260 168.260 42.490 168.290 ;
        RECT 42.830 168.260 43.060 168.290 ;
        RECT 43.310 169.040 43.690 169.260 ;
        RECT 43.310 168.260 43.540 169.040 ;
        RECT 43.880 168.590 44.110 169.260 ;
        RECT 44.360 168.940 44.640 169.260 ;
        RECT 44.360 168.590 44.590 168.940 ;
        RECT 43.880 168.260 44.590 168.590 ;
        RECT 41.990 168.090 42.280 168.100 ;
        RECT 41.940 167.790 42.340 168.090 ;
        RECT 44.090 167.840 44.390 168.260 ;
        RECT 45.190 167.540 45.590 170.240 ;
        RECT 46.840 169.390 47.240 169.690 ;
        RECT 46.940 167.640 47.140 169.390 ;
        RECT 34.640 166.440 46.040 167.540 ;
        RECT 46.840 167.340 47.240 167.640 ;
        RECT 39.640 165.940 41.340 166.440 ;
        RECT 47.420 165.980 48.070 180.830 ;
        RECT 70.220 180.240 70.670 180.280 ;
        RECT 48.640 179.990 50.745 180.240 ;
        RECT 68.635 179.990 70.740 180.240 ;
        RECT 48.720 179.410 50.570 179.990 ;
        RECT 70.220 179.930 70.670 179.990 ;
        RECT 72.020 179.680 72.170 180.830 ;
        RECT 72.320 179.680 72.550 180.380 ;
        RECT 72.020 179.530 72.550 179.680 ;
        RECT 48.640 179.160 50.745 179.410 ;
        RECT 68.635 179.380 70.740 179.410 ;
        RECT 72.320 179.380 72.550 179.530 ;
        RECT 72.760 179.830 72.990 180.380 ;
        RECT 73.170 180.230 73.570 180.530 ;
        RECT 75.135 180.405 75.425 180.450 ;
        RECT 76.115 180.405 76.405 180.450 ;
        RECT 77.095 180.405 77.385 180.450 ;
        RECT 78.075 180.405 78.365 180.450 ;
        RECT 80.195 180.430 80.485 180.450 ;
        RECT 81.175 180.430 81.465 180.450 ;
        RECT 82.155 180.430 82.445 180.450 ;
        RECT 83.135 180.430 83.425 180.450 ;
        RECT 80.170 180.405 83.520 180.430 ;
        RECT 75.135 180.255 78.970 180.405 ;
        RECT 73.320 179.830 73.470 180.230 ;
        RECT 75.135 180.220 75.425 180.255 ;
        RECT 76.115 180.220 76.405 180.255 ;
        RECT 77.095 180.220 77.385 180.255 ;
        RECT 78.075 180.220 78.365 180.255 ;
        RECT 72.760 179.680 73.470 179.830 ;
        RECT 72.760 179.380 72.990 179.680 ;
        RECT 66.720 179.180 70.740 179.380 ;
        RECT 48.640 178.530 50.745 178.580 ;
        RECT 48.640 178.330 54.370 178.530 ;
        RECT 48.640 177.500 50.745 177.750 ;
        RECT 48.920 176.920 50.220 177.500 ;
        RECT 48.640 176.670 50.745 176.920 ;
        RECT 48.640 175.840 50.745 176.090 ;
        RECT 48.870 175.260 50.170 175.840 ;
        RECT 48.640 175.010 50.745 175.260 ;
        RECT 48.640 174.180 50.745 174.430 ;
        RECT 48.970 173.600 50.270 174.180 ;
        RECT 51.770 173.980 52.170 174.280 ;
        RECT 48.640 173.350 50.745 173.600 ;
        RECT 48.640 172.655 50.745 172.770 ;
        RECT 48.220 172.520 50.745 172.655 ;
        RECT 48.220 172.505 49.095 172.520 ;
        RECT 48.220 170.930 48.370 172.505 ;
        RECT 48.640 171.930 50.745 171.940 ;
        RECT 51.870 171.930 52.020 173.980 ;
        RECT 48.640 171.780 52.020 171.930 ;
        RECT 48.640 171.690 50.745 171.780 ;
        RECT 48.220 170.630 48.620 170.930 ;
        RECT 51.870 169.180 52.020 171.780 ;
        RECT 54.170 170.430 54.370 178.330 ;
        RECT 54.070 170.130 54.470 170.430 ;
        RECT 60.020 170.180 60.420 179.030 ;
        RECT 48.710 168.950 53.070 169.180 ;
        RECT 48.720 168.930 53.070 168.950 ;
        RECT 48.500 167.080 48.730 168.790 ;
        RECT 48.980 168.230 49.210 168.790 ;
        RECT 48.870 167.930 49.270 168.230 ;
        RECT 48.420 166.780 48.820 167.080 ;
        RECT 48.980 166.790 49.210 167.930 ;
        RECT 49.460 167.080 49.690 168.790 ;
        RECT 49.940 168.230 50.170 168.790 ;
        RECT 49.870 167.930 50.270 168.230 ;
        RECT 49.370 166.780 49.770 167.080 ;
        RECT 49.940 166.790 50.170 167.930 ;
        RECT 50.420 167.080 50.650 168.790 ;
        RECT 50.320 166.780 50.720 167.080 ;
        RECT 51.120 166.630 51.320 168.930 ;
        RECT 51.560 168.780 51.790 168.790 ;
        RECT 51.470 168.480 51.870 168.780 ;
        RECT 51.560 166.790 51.790 168.480 ;
        RECT 52.040 167.630 52.270 168.790 ;
        RECT 52.520 168.780 52.750 168.790 ;
        RECT 52.420 168.480 52.820 168.780 ;
        RECT 51.970 167.330 52.370 167.630 ;
        RECT 52.040 166.790 52.270 167.330 ;
        RECT 52.520 166.790 52.750 168.480 ;
        RECT 53.000 167.630 53.230 168.790 ;
        RECT 53.480 168.780 53.710 168.790 ;
        RECT 53.420 168.480 53.820 168.780 ;
        RECT 52.920 167.330 53.320 167.630 ;
        RECT 53.000 166.790 53.230 167.330 ;
        RECT 53.480 166.790 53.710 168.480 ;
        RECT 54.170 167.630 54.370 170.130 ;
        RECT 54.870 169.630 60.970 170.180 ;
        RECT 54.795 169.055 59.845 169.305 ;
        RECT 54.070 167.330 54.470 167.630 ;
        RECT 54.795 166.630 55.045 169.055 ;
        RECT 55.520 169.040 55.810 169.055 ;
        RECT 56.480 169.040 56.770 169.055 ;
        RECT 58.580 169.040 58.870 169.055 ;
        RECT 59.540 169.040 59.830 169.055 ;
        RECT 55.220 168.580 55.620 168.880 ;
        RECT 55.310 166.835 55.540 168.580 ;
        RECT 55.790 168.230 56.020 168.835 ;
        RECT 56.170 168.580 56.570 168.880 ;
        RECT 55.720 167.930 56.120 168.230 ;
        RECT 55.790 166.835 56.020 167.930 ;
        RECT 56.270 166.835 56.500 168.580 ;
        RECT 56.750 168.230 56.980 168.835 ;
        RECT 57.120 168.580 57.520 168.880 ;
        RECT 56.670 167.930 57.070 168.230 ;
        RECT 56.750 166.835 56.980 167.930 ;
        RECT 57.230 166.835 57.460 168.580 ;
        RECT 58.370 167.080 58.600 168.835 ;
        RECT 58.850 167.630 59.080 168.835 ;
        RECT 58.770 167.330 59.170 167.630 ;
        RECT 58.270 166.780 58.670 167.080 ;
        RECT 58.850 166.835 59.080 167.330 ;
        RECT 59.330 167.080 59.560 168.835 ;
        RECT 59.810 167.630 60.040 168.835 ;
        RECT 59.720 167.330 60.120 167.630 ;
        RECT 59.270 166.780 59.670 167.080 ;
        RECT 59.810 166.835 60.040 167.330 ;
        RECT 60.290 167.080 60.520 168.835 ;
        RECT 61.270 168.530 61.670 173.130 ;
        RECT 66.720 171.380 66.920 179.180 ;
        RECT 68.635 179.160 70.740 179.180 ;
        RECT 72.510 179.105 72.800 179.175 ;
        RECT 71.920 178.955 72.800 179.105 ;
        RECT 67.370 178.580 67.770 178.880 ;
        RECT 67.495 171.405 67.645 178.580 ;
        RECT 68.635 178.330 70.740 178.580 ;
        RECT 69.070 177.750 70.370 178.330 ;
        RECT 68.635 177.500 70.740 177.750 ;
        RECT 68.635 176.670 70.740 176.920 ;
        RECT 70.970 176.730 71.370 177.030 ;
        RECT 69.020 176.090 70.320 176.670 ;
        RECT 68.635 175.840 70.740 176.090 ;
        RECT 68.635 175.010 70.740 175.260 ;
        RECT 68.920 174.430 70.220 175.010 ;
        RECT 68.635 174.180 70.740 174.430 ;
        RECT 71.070 174.280 71.220 176.730 ;
        RECT 71.370 176.230 71.770 176.530 ;
        RECT 70.920 173.980 71.320 174.280 ;
        RECT 68.635 173.350 70.740 173.600 ;
        RECT 69.020 172.770 70.320 173.350 ;
        RECT 70.970 172.780 71.370 173.080 ;
        RECT 68.635 172.520 70.740 172.770 ;
        RECT 71.020 171.980 71.320 172.780 ;
        RECT 68.635 171.690 70.740 171.940 ;
        RECT 70.270 171.680 70.570 171.690 ;
        RECT 70.970 171.680 71.370 171.980 ;
        RECT 66.620 171.080 67.020 171.380 ;
        RECT 67.495 171.255 69.920 171.405 ;
        RECT 67.870 170.180 68.170 170.580 ;
        RECT 68.470 170.530 68.770 170.930 ;
        RECT 60.220 166.780 60.620 167.080 ;
        RECT 61.820 166.780 62.220 169.980 ;
        RECT 62.370 168.180 62.770 169.430 ;
        RECT 63.810 169.030 64.100 169.080 ;
        RECT 63.620 168.830 64.120 169.030 ;
        RECT 64.720 168.830 65.120 169.130 ;
        RECT 63.620 168.690 63.770 168.830 ;
        RECT 67.170 168.780 67.570 169.080 ;
        RECT 63.600 167.930 63.830 168.690 ;
        RECT 64.080 168.480 64.310 168.690 ;
        RECT 63.970 168.180 64.370 168.480 ;
        RECT 63.520 167.630 63.920 167.930 ;
        RECT 49.170 166.380 53.520 166.630 ;
        RECT 54.795 166.380 60.345 166.630 ;
        RECT 39.590 164.240 41.390 165.940 ;
        RECT 47.420 165.580 54.220 165.980 ;
        RECT 57.770 165.580 58.120 166.380 ;
        RECT 62.370 166.130 62.770 167.330 ;
        RECT 63.600 166.790 63.830 167.630 ;
        RECT 64.080 166.790 64.310 168.180 ;
        RECT 64.560 167.930 64.790 168.690 ;
        RECT 64.470 167.630 64.870 167.930 ;
        RECT 64.560 166.790 64.790 167.630 ;
        RECT 65.040 167.330 65.270 168.690 ;
        RECT 65.520 167.930 65.750 168.690 ;
        RECT 65.420 167.630 65.820 167.930 ;
        RECT 64.970 167.030 65.370 167.330 ;
        RECT 65.040 166.790 65.270 167.030 ;
        RECT 65.520 166.790 65.750 167.630 ;
        RECT 66.470 166.630 66.870 167.930 ;
        RECT 67.320 167.830 67.470 168.780 ;
        RECT 67.170 167.530 67.570 167.830 ;
        RECT 67.320 166.630 67.470 167.530 ;
        RECT 64.220 166.330 64.620 166.630 ;
        RECT 65.220 166.380 66.870 166.630 ;
        RECT 66.470 165.980 66.870 166.380 ;
        RECT 67.170 166.330 67.570 166.630 ;
        RECT 67.920 166.455 68.070 170.180 ;
        RECT 68.520 166.855 68.670 170.530 ;
        RECT 68.870 167.530 69.270 167.830 ;
        RECT 69.770 167.530 69.920 171.255 ;
        RECT 70.420 170.730 70.570 171.680 ;
        RECT 70.320 170.430 70.720 170.730 ;
        RECT 70.470 167.530 70.870 167.830 ;
        RECT 68.970 167.030 69.200 167.530 ;
        RECT 69.760 167.030 69.990 167.530 ;
        RECT 70.550 167.030 70.780 167.530 ;
        RECT 69.250 166.855 69.710 166.870 ;
        RECT 68.520 166.705 69.710 166.855 ;
        RECT 69.250 166.640 69.710 166.705 ;
        RECT 70.040 166.640 70.500 166.870 ;
        RECT 70.195 166.455 70.345 166.640 ;
        RECT 67.920 166.305 70.345 166.455 ;
        RECT 71.620 165.980 71.770 176.230 ;
        RECT 71.920 175.130 72.070 178.955 ;
        RECT 72.510 178.945 72.800 178.955 ;
        RECT 72.510 177.430 72.800 177.440 ;
        RECT 72.470 177.230 73.420 177.430 ;
        RECT 72.510 177.210 72.800 177.230 ;
        RECT 72.320 177.030 72.550 177.050 ;
        RECT 72.220 176.730 72.620 177.030 ;
        RECT 72.320 176.050 72.550 176.730 ;
        RECT 72.760 176.530 72.990 177.050 ;
        RECT 72.720 176.230 73.120 176.530 ;
        RECT 72.760 176.050 72.990 176.230 ;
        RECT 72.510 175.130 72.800 175.180 ;
        RECT 71.920 174.980 72.820 175.130 ;
        RECT 71.920 166.555 72.070 174.980 ;
        RECT 72.510 174.950 72.800 174.980 ;
        RECT 72.320 171.380 72.550 174.790 ;
        RECT 72.220 171.080 72.620 171.380 ;
        RECT 72.320 166.790 72.550 171.080 ;
        RECT 72.760 167.130 72.990 174.790 ;
        RECT 73.270 168.030 73.420 177.230 ;
        RECT 73.570 176.480 73.970 176.780 ;
        RECT 73.570 169.980 73.720 176.480 ;
        RECT 73.870 175.530 74.270 175.830 ;
        RECT 73.970 171.980 74.170 175.530 ;
        RECT 74.430 174.930 74.660 180.015 ;
        RECT 74.920 176.780 75.150 180.015 ;
        RECT 74.820 176.480 75.220 176.780 ;
        RECT 74.320 174.630 74.720 174.930 ;
        RECT 74.430 174.015 74.660 174.630 ;
        RECT 74.920 174.015 75.150 176.480 ;
        RECT 75.410 174.930 75.640 180.015 ;
        RECT 75.900 176.780 76.130 180.015 ;
        RECT 75.820 176.480 76.220 176.780 ;
        RECT 75.320 174.630 75.720 174.930 ;
        RECT 75.410 174.015 75.640 174.630 ;
        RECT 75.900 174.015 76.130 176.480 ;
        RECT 76.390 174.930 76.620 180.015 ;
        RECT 76.880 176.780 77.110 180.015 ;
        RECT 76.820 176.480 77.220 176.780 ;
        RECT 76.270 174.630 76.670 174.930 ;
        RECT 76.390 174.015 76.620 174.630 ;
        RECT 76.880 174.015 77.110 176.480 ;
        RECT 77.370 174.930 77.600 180.015 ;
        RECT 77.860 176.780 78.090 180.015 ;
        RECT 77.770 176.480 78.170 176.780 ;
        RECT 77.270 174.630 77.670 174.930 ;
        RECT 77.370 174.015 77.600 174.630 ;
        RECT 77.860 174.015 78.090 176.480 ;
        RECT 78.350 174.930 78.580 180.015 ;
        RECT 78.820 177.630 78.970 180.255 ;
        RECT 80.170 180.255 84.020 180.405 ;
        RECT 80.170 180.230 83.520 180.255 ;
        RECT 80.195 180.220 80.485 180.230 ;
        RECT 81.175 180.220 81.465 180.230 ;
        RECT 82.155 180.220 82.445 180.230 ;
        RECT 83.135 180.220 83.425 180.230 ;
        RECT 78.720 177.330 79.120 177.630 ;
        RECT 78.270 174.630 78.670 174.930 ;
        RECT 78.350 174.015 78.580 174.630 ;
        RECT 74.645 173.755 74.935 173.810 ;
        RECT 75.625 173.755 75.915 173.810 ;
        RECT 76.605 173.755 76.895 173.810 ;
        RECT 77.585 173.755 77.875 173.810 ;
        RECT 78.820 173.755 78.970 177.330 ;
        RECT 79.490 174.930 79.720 180.015 ;
        RECT 79.980 175.830 80.210 180.015 ;
        RECT 79.870 175.530 80.270 175.830 ;
        RECT 79.420 174.630 79.820 174.930 ;
        RECT 79.490 174.015 79.720 174.630 ;
        RECT 79.980 174.015 80.210 175.530 ;
        RECT 80.470 174.930 80.700 180.015 ;
        RECT 80.960 175.830 81.190 180.015 ;
        RECT 80.870 175.530 81.270 175.830 ;
        RECT 80.370 174.630 80.770 174.930 ;
        RECT 80.470 174.015 80.700 174.630 ;
        RECT 80.960 174.015 81.190 175.530 ;
        RECT 81.450 174.930 81.680 180.015 ;
        RECT 81.940 175.830 82.170 180.015 ;
        RECT 81.870 175.530 82.270 175.830 ;
        RECT 81.370 174.630 81.770 174.930 ;
        RECT 81.450 174.015 81.680 174.630 ;
        RECT 81.940 174.015 82.170 175.530 ;
        RECT 82.430 174.930 82.660 180.015 ;
        RECT 82.920 175.830 83.150 180.015 ;
        RECT 82.820 175.530 83.220 175.830 ;
        RECT 82.370 174.630 82.770 174.930 ;
        RECT 82.430 174.015 82.660 174.630 ;
        RECT 82.920 174.015 83.150 175.530 ;
        RECT 83.410 174.930 83.640 180.015 ;
        RECT 83.870 178.230 84.020 180.255 ;
        RECT 84.170 178.880 84.370 180.830 ;
        RECT 84.770 180.180 101.670 180.580 ;
        RECT 92.720 180.015 92.920 180.180 ;
        RECT 84.540 178.880 84.770 180.015 ;
        RECT 85.330 178.880 85.560 180.015 ;
        RECT 84.170 178.630 85.560 178.880 ;
        RECT 83.820 177.930 84.220 178.230 ;
        RECT 83.320 174.630 83.720 174.930 ;
        RECT 83.410 174.015 83.640 174.630 ;
        RECT 79.670 173.755 80.070 173.830 ;
        RECT 80.685 173.755 80.975 173.810 ;
        RECT 81.665 173.755 81.955 173.810 ;
        RECT 82.645 173.755 82.935 173.810 ;
        RECT 83.870 173.755 84.020 177.930 ;
        RECT 74.645 173.605 79.345 173.755 ;
        RECT 74.645 173.580 74.935 173.605 ;
        RECT 75.625 173.580 75.915 173.605 ;
        RECT 76.605 173.580 76.895 173.605 ;
        RECT 77.585 173.580 77.875 173.605 ;
        RECT 74.645 173.255 74.935 173.270 ;
        RECT 75.625 173.255 75.915 173.270 ;
        RECT 76.605 173.255 76.895 173.270 ;
        RECT 77.585 173.255 77.875 173.270 ;
        RECT 78.270 173.255 78.670 173.380 ;
        RECT 79.195 173.255 79.345 173.605 ;
        RECT 79.670 173.605 84.020 173.755 ;
        RECT 79.670 173.530 80.070 173.605 ;
        RECT 80.685 173.580 80.975 173.605 ;
        RECT 81.665 173.580 81.955 173.605 ;
        RECT 82.645 173.580 82.935 173.605 ;
        RECT 79.705 173.255 79.995 173.270 ;
        RECT 80.685 173.255 80.975 173.270 ;
        RECT 81.665 173.255 81.955 173.270 ;
        RECT 82.645 173.255 82.935 173.270 ;
        RECT 74.645 173.105 78.970 173.255 ;
        RECT 79.195 173.105 84.020 173.255 ;
        RECT 74.645 173.040 74.935 173.105 ;
        RECT 75.625 173.040 75.915 173.105 ;
        RECT 76.605 173.040 76.895 173.105 ;
        RECT 77.585 173.040 77.875 173.105 ;
        RECT 78.270 173.080 78.670 173.105 ;
        RECT 74.430 172.630 74.660 172.835 ;
        RECT 74.320 172.330 74.720 172.630 ;
        RECT 73.870 171.680 74.270 171.980 ;
        RECT 73.570 169.680 73.970 169.980 ;
        RECT 73.170 167.730 73.570 168.030 ;
        RECT 72.760 166.880 73.520 167.130 ;
        RECT 72.760 166.790 72.990 166.880 ;
        RECT 72.470 166.555 72.870 166.630 ;
        RECT 71.920 166.405 72.870 166.555 ;
        RECT 72.470 166.330 72.870 166.405 ;
        RECT 73.220 165.980 73.520 166.880 ;
        RECT 74.430 166.835 74.660 172.330 ;
        RECT 74.920 171.980 75.150 172.835 ;
        RECT 75.410 172.630 75.640 172.835 ;
        RECT 75.320 172.330 75.720 172.630 ;
        RECT 74.820 171.680 75.220 171.980 ;
        RECT 74.920 166.835 75.150 171.680 ;
        RECT 75.410 166.835 75.640 172.330 ;
        RECT 75.900 171.980 76.130 172.835 ;
        RECT 76.390 172.630 76.620 172.835 ;
        RECT 76.270 172.330 76.670 172.630 ;
        RECT 75.820 171.680 76.220 171.980 ;
        RECT 75.900 166.835 76.130 171.680 ;
        RECT 76.390 166.835 76.620 172.330 ;
        RECT 76.880 171.980 77.110 172.835 ;
        RECT 77.370 172.630 77.600 172.835 ;
        RECT 77.270 172.330 77.670 172.630 ;
        RECT 76.820 171.680 77.220 171.980 ;
        RECT 76.880 166.835 77.110 171.680 ;
        RECT 77.370 166.835 77.600 172.330 ;
        RECT 77.860 171.980 78.090 172.835 ;
        RECT 78.350 172.630 78.580 172.835 ;
        RECT 78.270 172.330 78.670 172.630 ;
        RECT 77.770 171.680 78.170 171.980 ;
        RECT 77.860 166.835 78.090 171.680 ;
        RECT 78.350 166.835 78.580 172.330 ;
        RECT 75.135 166.605 75.425 166.630 ;
        RECT 76.115 166.605 76.405 166.630 ;
        RECT 77.095 166.605 77.385 166.630 ;
        RECT 78.075 166.605 78.365 166.630 ;
        RECT 78.820 166.605 78.970 173.105 ;
        RECT 79.705 173.040 79.995 173.105 ;
        RECT 80.685 173.040 80.975 173.105 ;
        RECT 81.665 173.040 81.955 173.105 ;
        RECT 82.645 173.040 82.935 173.105 ;
        RECT 79.490 172.630 79.720 172.835 ;
        RECT 79.420 172.330 79.820 172.630 ;
        RECT 79.490 166.835 79.720 172.330 ;
        RECT 79.980 169.980 80.210 172.835 ;
        RECT 80.470 172.630 80.700 172.835 ;
        RECT 80.370 172.330 80.770 172.630 ;
        RECT 79.870 169.680 80.270 169.980 ;
        RECT 79.980 166.835 80.210 169.680 ;
        RECT 80.470 166.835 80.700 172.330 ;
        RECT 80.960 169.980 81.190 172.835 ;
        RECT 81.450 172.630 81.680 172.835 ;
        RECT 81.370 172.330 81.770 172.630 ;
        RECT 80.870 169.680 81.270 169.980 ;
        RECT 80.960 166.835 81.190 169.680 ;
        RECT 81.450 166.835 81.680 172.330 ;
        RECT 81.940 169.980 82.170 172.835 ;
        RECT 82.430 172.630 82.660 172.835 ;
        RECT 82.320 172.330 82.720 172.630 ;
        RECT 81.870 169.680 82.270 169.980 ;
        RECT 81.940 166.835 82.170 169.680 ;
        RECT 82.430 166.835 82.660 172.330 ;
        RECT 82.920 169.980 83.150 172.835 ;
        RECT 83.410 172.630 83.640 172.835 ;
        RECT 83.320 172.330 83.720 172.630 ;
        RECT 82.820 169.680 83.220 169.980 ;
        RECT 82.920 166.835 83.150 169.680 ;
        RECT 83.410 166.835 83.640 172.330 ;
        RECT 75.135 166.455 78.970 166.605 ;
        RECT 80.195 166.605 80.485 166.630 ;
        RECT 81.175 166.605 81.465 166.630 ;
        RECT 82.155 166.605 82.445 166.630 ;
        RECT 83.135 166.605 83.425 166.630 ;
        RECT 83.870 166.605 84.020 173.105 ;
        RECT 84.540 172.015 84.770 178.630 ;
        RECT 85.330 172.015 85.560 178.630 ;
        RECT 85.900 175.730 86.130 180.015 ;
        RECT 86.690 178.980 86.920 180.015 ;
        RECT 86.620 178.680 87.020 178.980 ;
        RECT 86.690 176.490 86.920 178.680 ;
        RECT 86.640 176.190 87.040 176.490 ;
        RECT 85.820 175.430 86.220 175.730 ;
        RECT 85.900 172.015 86.130 175.430 ;
        RECT 86.690 173.440 86.920 176.190 ;
        RECT 87.260 174.290 87.490 180.015 ;
        RECT 88.050 178.980 88.280 180.015 ;
        RECT 87.970 178.680 88.370 178.980 ;
        RECT 88.050 176.490 88.280 178.680 ;
        RECT 87.990 176.190 88.390 176.490 ;
        RECT 87.190 173.990 87.590 174.290 ;
        RECT 86.640 173.140 87.040 173.440 ;
        RECT 86.690 172.015 86.920 173.140 ;
        RECT 87.260 172.015 87.490 173.990 ;
        RECT 88.050 173.440 88.280 176.190 ;
        RECT 88.620 174.890 88.850 180.015 ;
        RECT 89.410 178.980 89.640 180.015 ;
        RECT 89.320 178.680 89.720 178.980 ;
        RECT 89.410 176.490 89.640 178.680 ;
        RECT 89.340 176.190 89.740 176.490 ;
        RECT 88.540 174.590 88.940 174.890 ;
        RECT 87.990 173.140 88.390 173.440 ;
        RECT 88.050 172.015 88.280 173.140 ;
        RECT 88.620 172.650 88.850 174.590 ;
        RECT 89.410 173.440 89.640 176.190 ;
        RECT 89.980 174.890 90.210 180.015 ;
        RECT 90.770 178.980 91.000 180.015 ;
        RECT 90.670 178.680 91.070 178.980 ;
        RECT 90.770 176.490 91.000 178.680 ;
        RECT 90.690 176.190 91.090 176.490 ;
        RECT 89.890 174.590 90.290 174.890 ;
        RECT 89.340 173.140 89.740 173.440 ;
        RECT 88.560 172.350 88.960 172.650 ;
        RECT 88.620 172.015 88.850 172.350 ;
        RECT 89.410 172.015 89.640 173.140 ;
        RECT 89.980 172.650 90.210 174.590 ;
        RECT 90.770 173.440 91.000 176.190 ;
        RECT 91.340 174.890 91.570 180.015 ;
        RECT 92.130 178.980 92.360 180.015 ;
        RECT 92.070 178.680 92.470 178.980 ;
        RECT 92.130 176.490 92.360 178.680 ;
        RECT 92.090 176.190 92.490 176.490 ;
        RECT 91.290 174.590 91.690 174.890 ;
        RECT 90.690 173.140 91.090 173.440 ;
        RECT 89.910 172.350 90.310 172.650 ;
        RECT 89.980 172.015 90.210 172.350 ;
        RECT 90.770 172.015 91.000 173.140 ;
        RECT 91.340 172.650 91.570 174.590 ;
        RECT 92.130 173.440 92.360 176.190 ;
        RECT 92.090 173.140 92.490 173.440 ;
        RECT 91.310 172.350 91.710 172.650 ;
        RECT 91.340 172.015 91.570 172.350 ;
        RECT 92.130 172.015 92.360 173.140 ;
        RECT 92.700 172.015 92.930 180.015 ;
        RECT 93.490 178.980 93.720 180.015 ;
        RECT 93.420 178.680 93.820 178.980 ;
        RECT 93.490 176.490 93.720 178.680 ;
        RECT 93.440 176.190 93.840 176.490 ;
        RECT 93.490 173.440 93.720 176.190 ;
        RECT 94.060 174.890 94.290 180.015 ;
        RECT 94.850 178.980 95.080 180.015 ;
        RECT 94.770 178.680 95.170 178.980 ;
        RECT 94.850 176.490 95.080 178.680 ;
        RECT 94.790 176.190 95.190 176.490 ;
        RECT 93.990 174.590 94.390 174.890 ;
        RECT 93.440 173.140 93.840 173.440 ;
        RECT 93.490 172.015 93.720 173.140 ;
        RECT 94.060 172.650 94.290 174.590 ;
        RECT 94.850 173.440 95.080 176.190 ;
        RECT 95.420 174.890 95.650 180.015 ;
        RECT 96.210 178.980 96.440 180.015 ;
        RECT 96.120 178.680 96.520 178.980 ;
        RECT 96.210 176.490 96.440 178.680 ;
        RECT 96.140 176.190 96.540 176.490 ;
        RECT 95.340 174.590 95.740 174.890 ;
        RECT 94.790 173.140 95.190 173.440 ;
        RECT 94.010 172.350 94.410 172.650 ;
        RECT 94.060 172.015 94.290 172.350 ;
        RECT 94.850 172.015 95.080 173.140 ;
        RECT 95.420 172.650 95.650 174.590 ;
        RECT 96.210 173.440 96.440 176.190 ;
        RECT 96.780 174.890 97.010 180.015 ;
        RECT 97.570 178.980 97.800 180.015 ;
        RECT 97.470 178.680 97.870 178.980 ;
        RECT 97.570 176.490 97.800 178.680 ;
        RECT 97.490 176.190 97.890 176.490 ;
        RECT 96.690 174.590 97.090 174.890 ;
        RECT 96.140 173.140 96.540 173.440 ;
        RECT 95.360 172.350 95.760 172.650 ;
        RECT 95.420 172.015 95.650 172.350 ;
        RECT 96.210 172.015 96.440 173.140 ;
        RECT 96.780 172.650 97.010 174.590 ;
        RECT 97.570 173.440 97.800 176.190 ;
        RECT 98.140 175.740 98.370 180.015 ;
        RECT 98.930 178.980 99.160 180.015 ;
        RECT 98.870 178.680 99.270 178.980 ;
        RECT 98.930 176.490 99.160 178.680 ;
        RECT 98.890 176.190 99.290 176.490 ;
        RECT 98.090 175.440 98.490 175.740 ;
        RECT 97.490 173.140 97.890 173.440 ;
        RECT 96.710 172.350 97.110 172.650 ;
        RECT 96.780 172.015 97.010 172.350 ;
        RECT 97.570 172.015 97.800 173.140 ;
        RECT 98.140 172.015 98.370 175.440 ;
        RECT 98.930 173.440 99.160 176.190 ;
        RECT 99.500 175.740 99.730 180.015 ;
        RECT 100.290 178.980 100.520 180.015 ;
        RECT 100.860 178.980 101.090 180.015 ;
        RECT 101.650 178.980 101.880 180.015 ;
        RECT 102.320 178.980 102.970 180.830 ;
        RECT 100.220 178.680 100.620 178.980 ;
        RECT 100.860 178.730 102.970 178.980 ;
        RECT 100.290 176.490 100.520 178.680 ;
        RECT 100.240 176.190 100.640 176.490 ;
        RECT 99.440 175.440 99.840 175.740 ;
        RECT 98.890 173.140 99.290 173.440 ;
        RECT 98.930 172.015 99.160 173.140 ;
        RECT 99.500 172.015 99.730 175.440 ;
        RECT 100.290 173.440 100.520 176.190 ;
        RECT 100.240 173.140 100.640 173.440 ;
        RECT 100.290 172.015 100.520 173.140 ;
        RECT 100.860 172.015 101.090 178.730 ;
        RECT 101.650 172.015 101.880 178.730 ;
        RECT 92.720 171.830 92.920 172.015 ;
        RECT 84.770 171.430 101.670 171.830 ;
        RECT 102.320 171.180 102.970 178.730 ;
        RECT 103.120 175.430 103.520 175.730 ;
        RECT 86.420 170.480 86.820 170.780 ;
        RECT 86.470 170.140 86.720 170.480 ;
        RECT 92.450 170.180 92.680 170.710 ;
        RECT 93.740 170.180 93.970 170.710 ;
        RECT 95.030 170.230 95.260 170.710 ;
        RECT 95.670 170.530 102.970 171.180 ;
        RECT 86.470 170.130 86.760 170.140 ;
        RECT 88.570 170.130 88.860 170.140 ;
        RECT 86.470 169.930 88.870 170.130 ;
        RECT 86.470 169.910 86.760 169.930 ;
        RECT 87.320 169.750 87.520 169.930 ;
        RECT 88.570 169.910 88.860 169.930 ;
        RECT 92.370 169.880 92.770 170.180 ;
        RECT 93.670 169.880 94.070 170.180 ;
        RECT 95.030 170.080 95.570 170.230 ;
        RECT 103.220 170.180 103.420 175.430 ;
        RECT 85.210 168.930 85.440 169.750 ;
        RECT 85.690 168.930 85.920 169.750 ;
        RECT 86.260 169.030 86.490 169.750 ;
        RECT 85.210 168.780 85.920 168.930 ;
        RECT 85.210 168.530 85.440 168.780 ;
        RECT 85.690 168.580 85.920 168.780 ;
        RECT 86.170 168.730 86.570 169.030 ;
        RECT 85.620 168.530 86.020 168.580 ;
        RECT 85.210 168.330 86.020 168.530 ;
        RECT 85.210 167.750 85.440 168.330 ;
        RECT 85.620 168.280 86.020 168.330 ;
        RECT 85.690 167.750 85.920 168.280 ;
        RECT 86.260 167.750 86.490 168.730 ;
        RECT 86.740 168.580 86.970 169.750 ;
        RECT 86.670 168.280 87.070 168.580 ;
        RECT 86.740 167.750 86.970 168.280 ;
        RECT 87.310 167.750 87.540 169.750 ;
        RECT 87.790 168.580 88.020 169.750 ;
        RECT 88.360 169.030 88.590 169.750 ;
        RECT 88.270 168.730 88.670 169.030 ;
        RECT 87.720 168.280 88.120 168.580 ;
        RECT 87.790 167.750 88.020 168.280 ;
        RECT 88.360 167.750 88.590 168.730 ;
        RECT 88.840 168.580 89.070 169.750 ;
        RECT 89.410 168.980 89.640 169.750 ;
        RECT 89.890 168.980 90.120 169.750 ;
        RECT 92.450 169.710 92.680 169.880 ;
        RECT 93.740 169.710 93.970 169.880 ;
        RECT 95.030 169.710 95.260 170.080 ;
        RECT 92.730 169.275 93.690 169.505 ;
        RECT 94.020 169.275 94.980 169.505 ;
        RECT 89.410 168.830 90.120 168.980 ;
        RECT 88.770 168.280 89.170 168.580 ;
        RECT 89.410 168.530 89.640 168.830 ;
        RECT 89.890 168.580 90.120 168.830 ;
        RECT 89.820 168.530 90.220 168.580 ;
        RECT 93.120 168.530 93.320 169.275 ;
        RECT 94.420 168.980 94.620 169.275 ;
        RECT 94.320 168.680 94.720 168.980 ;
        RECT 89.410 168.330 90.670 168.530 ;
        RECT 88.840 167.750 89.070 168.280 ;
        RECT 89.410 167.750 89.640 168.330 ;
        RECT 89.820 168.280 90.220 168.330 ;
        RECT 89.890 167.750 90.120 168.280 ;
        RECT 87.320 167.590 87.520 167.750 ;
        RECT 85.420 167.580 85.710 167.590 ;
        RECT 87.320 167.580 87.810 167.590 ;
        RECT 89.620 167.580 89.910 167.590 ;
        RECT 85.320 167.380 89.970 167.580 ;
        RECT 85.420 167.360 85.710 167.380 ;
        RECT 87.520 167.360 87.810 167.380 ;
        RECT 89.620 167.360 89.910 167.380 ;
        RECT 80.195 166.455 84.020 166.605 ;
        RECT 75.135 166.400 75.425 166.455 ;
        RECT 76.115 166.400 76.405 166.455 ;
        RECT 77.095 166.400 77.385 166.455 ;
        RECT 78.075 166.400 78.365 166.455 ;
        RECT 80.195 166.400 80.485 166.455 ;
        RECT 81.175 166.400 81.465 166.455 ;
        RECT 82.155 166.400 82.445 166.455 ;
        RECT 83.135 166.400 83.425 166.455 ;
        RECT 90.420 165.980 90.670 168.330 ;
        RECT 93.020 168.230 93.420 168.530 ;
        RECT 95.420 167.330 95.570 170.080 ;
        RECT 103.120 169.880 103.520 170.180 ;
        RECT 101.360 169.780 101.730 169.860 ;
        RECT 100.470 169.630 101.730 169.780 ;
        RECT 98.820 169.080 99.220 169.380 ;
        RECT 95.220 167.030 95.620 167.330 ;
        RECT 98.920 166.680 99.120 169.080 ;
        RECT 100.470 168.030 100.620 169.630 ;
        RECT 101.360 169.550 101.730 169.630 ;
        RECT 101.760 169.380 102.150 169.395 ;
        RECT 103.990 169.390 104.140 169.440 ;
        RECT 101.760 169.095 102.170 169.380 ;
        RECT 101.770 169.080 102.170 169.095 ;
        RECT 103.840 169.315 104.240 169.390 ;
        RECT 105.440 169.315 105.590 184.490 ;
        RECT 103.840 169.165 105.590 169.315 ;
        RECT 103.840 169.090 104.240 169.165 ;
        RECT 101.040 168.280 102.420 168.290 ;
        RECT 100.370 167.730 100.770 168.030 ;
        RECT 98.820 166.380 99.220 166.680 ;
        RECT 100.920 165.980 102.970 168.280 ;
        RECT 63.120 165.580 73.520 165.980 ;
        RECT 84.720 165.580 102.970 165.980 ;
        RECT 47.420 164.880 102.970 165.580 ;
        RECT 66.840 164.240 68.640 164.880 ;
        RECT 105.190 163.865 105.590 163.990 ;
        RECT 32.590 163.715 105.590 163.865 ;
        RECT 105.190 163.690 105.590 163.715 ;
        RECT 105.840 163.540 105.990 185.115 ;
        RECT 80.315 163.390 105.990 163.540 ;
        RECT 32.265 163.090 80.015 163.240 ;
        RECT 80.315 163.140 80.615 163.390 ;
        RECT 106.140 163.240 106.290 185.565 ;
        RECT 31.965 162.790 79.565 162.940 ;
        RECT 79.715 162.840 80.015 163.090 ;
        RECT 80.765 163.090 106.290 163.240 ;
        RECT 80.765 162.840 81.065 163.090 ;
        RECT 106.440 162.940 106.590 186.015 ;
        RECT 31.665 162.490 79.115 162.640 ;
        RECT 79.265 162.540 79.565 162.790 ;
        RECT 81.215 162.790 106.590 162.940 ;
        RECT 81.215 162.540 81.515 162.790 ;
        RECT 106.740 162.640 106.890 186.315 ;
        RECT 31.365 162.190 78.665 162.340 ;
        RECT 78.815 162.240 79.115 162.490 ;
        RECT 81.665 162.490 106.890 162.640 ;
        RECT 81.665 162.240 81.965 162.490 ;
        RECT 107.040 162.340 107.190 187.515 ;
        RECT 110.490 187.490 110.890 187.515 ;
        RECT 119.690 187.315 120.090 187.440 ;
        RECT 31.065 161.890 78.215 162.040 ;
        RECT 78.365 161.940 78.665 162.190 ;
        RECT 82.115 162.190 107.190 162.340 ;
        RECT 107.340 187.165 120.090 187.315 ;
        RECT 82.115 161.940 82.415 162.190 ;
        RECT 107.340 162.040 107.490 187.165 ;
        RECT 119.690 187.140 120.090 187.165 ;
        RECT 133.490 186.965 133.890 187.090 ;
        RECT 30.765 161.590 77.765 161.740 ;
        RECT 77.915 161.640 78.215 161.890 ;
        RECT 82.565 161.890 107.490 162.040 ;
        RECT 107.640 186.815 133.890 186.965 ;
        RECT 82.565 161.640 82.865 161.890 ;
        RECT 107.640 161.740 107.790 186.815 ;
        RECT 133.490 186.790 133.890 186.815 ;
        RECT 128.890 186.515 129.290 186.640 ;
        RECT 107.940 186.365 129.290 186.515 ;
        RECT 107.940 183.590 108.090 186.365 ;
        RECT 128.890 186.340 129.290 186.365 ;
        RECT 142.690 186.590 143.090 186.640 ;
        RECT 145.790 186.590 146.190 186.640 ;
        RECT 142.690 186.440 146.190 186.590 ;
        RECT 142.690 186.340 143.090 186.440 ;
        RECT 145.790 186.340 146.190 186.440 ;
        RECT 147.990 186.190 148.390 186.340 ;
        RECT 108.415 186.040 148.390 186.190 ;
        RECT 107.940 183.190 108.240 183.590 ;
        RECT 108.415 183.140 108.565 186.040 ;
        RECT 150.070 185.865 150.210 219.940 ;
        RECT 150.600 219.290 150.900 219.690 ;
        RECT 108.790 185.715 150.215 185.865 ;
        RECT 108.790 184.840 108.940 185.715 ;
        RECT 109.245 185.065 141.595 185.515 ;
        RECT 141.795 185.065 149.245 185.515 ;
        RECT 108.740 184.440 109.040 184.840 ;
        RECT 108.390 182.740 108.690 183.140 ;
        RECT 109.245 180.215 109.745 185.065 ;
        RECT 115.190 185.040 117.140 185.065 ;
        RECT 141.395 184.775 141.595 185.065 ;
        RECT 125.145 184.715 125.545 184.765 ;
        RECT 110.245 184.465 140.845 184.715 ;
        RECT 109.965 180.215 110.195 184.270 ;
        RECT 120.255 180.215 120.485 184.270 ;
        RECT 130.545 180.215 130.775 184.270 ;
        RECT 140.835 180.215 141.065 184.270 ;
        RECT 141.365 182.415 141.625 184.775 ;
        RECT 141.815 184.690 145.090 185.065 ;
        RECT 141.815 184.660 144.575 184.690 ;
        RECT 145.740 184.490 146.140 184.790 ;
        RECT 147.390 184.715 147.790 184.790 ;
        RECT 147.390 184.490 147.795 184.715 ;
        RECT 147.990 184.490 148.390 184.790 ;
        RECT 145.890 183.915 146.040 184.490 ;
        RECT 144.095 183.875 144.545 183.915 ;
        RECT 143.295 183.855 143.695 183.865 ;
        RECT 142.485 183.555 142.935 183.855 ;
        RECT 143.240 183.565 143.695 183.855 ;
        RECT 144.085 183.565 144.545 183.875 ;
        RECT 145.745 183.615 146.145 183.915 ;
        RECT 142.115 183.365 142.425 183.425 ;
        RECT 141.995 183.065 142.425 183.365 ;
        RECT 142.115 183.005 142.425 183.065 ;
        RECT 142.635 182.975 142.795 183.555 ;
        RECT 143.240 183.545 143.690 183.565 ;
        RECT 144.085 183.545 144.540 183.565 ;
        RECT 143.715 183.015 144.025 183.125 ;
        RECT 143.645 182.975 144.045 183.015 ;
        RECT 142.635 182.750 144.045 182.975 ;
        RECT 143.645 182.715 144.045 182.750 ;
        RECT 143.715 182.705 144.025 182.715 ;
        RECT 141.815 182.415 144.575 182.420 ;
        RECT 141.365 181.965 144.575 182.415 ;
        RECT 141.365 180.215 141.625 181.965 ;
        RECT 141.815 181.940 144.575 181.965 ;
        RECT 142.095 181.680 142.495 181.700 ;
        RECT 142.085 181.400 142.495 181.680 ;
        RECT 142.085 181.370 142.455 181.400 ;
        RECT 145.895 180.815 146.045 183.615 ;
        RECT 146.245 183.165 146.645 183.465 ;
        RECT 142.495 180.505 142.920 180.810 ;
        RECT 143.240 180.505 143.695 180.815 ;
        RECT 109.245 178.515 141.625 180.215 ;
        RECT 142.695 180.165 142.845 180.505 ;
        RECT 144.085 180.485 144.545 180.815 ;
        RECT 145.745 180.515 146.145 180.815 ;
        RECT 144.095 180.465 144.545 180.485 ;
        RECT 143.295 180.235 143.695 180.265 ;
        RECT 143.280 180.165 143.705 180.235 ;
        RECT 142.695 180.015 143.705 180.165 ;
        RECT 143.280 179.930 143.705 180.015 ;
        RECT 145.345 179.965 145.745 180.265 ;
        RECT 141.815 179.220 145.035 179.700 ;
        RECT 143.730 179.015 144.140 179.070 ;
        RECT 143.730 178.965 144.195 179.015 ;
        RECT 142.085 178.585 142.505 178.945 ;
        RECT 142.745 178.815 144.195 178.965 ;
        RECT 108.640 173.760 109.040 174.060 ;
        RECT 108.190 169.310 108.590 169.610 ;
        RECT 108.340 168.690 108.490 169.310 ;
        RECT 108.190 168.390 108.590 168.690 ;
        RECT 108.790 168.040 108.940 173.760 ;
        RECT 108.540 167.740 108.940 168.040 ;
        RECT 109.245 168.015 109.745 178.515 ;
        RECT 109.965 174.270 110.195 178.515 ;
        RECT 120.255 174.270 120.485 178.515 ;
        RECT 130.545 174.270 130.775 178.515 ;
        RECT 140.835 174.270 141.065 178.515 ;
        RECT 141.365 176.965 141.625 178.515 ;
        RECT 142.745 178.415 142.895 178.815 ;
        RECT 143.795 178.715 144.195 178.815 ;
        RECT 143.250 178.515 143.625 178.525 ;
        RECT 142.485 178.115 142.935 178.415 ;
        RECT 143.195 177.715 143.645 178.515 ;
        RECT 143.785 178.135 144.205 178.495 ;
        RECT 144.715 178.465 145.145 178.575 ;
        RECT 144.695 178.165 145.145 178.465 ;
        RECT 143.945 177.465 144.095 178.135 ;
        RECT 144.715 178.105 145.145 178.165 ;
        RECT 144.795 178.100 145.145 178.105 ;
        RECT 144.795 177.515 144.995 178.100 ;
        RECT 143.445 177.215 144.095 177.465 ;
        RECT 144.695 177.215 145.095 177.515 ;
        RECT 143.445 177.165 143.845 177.215 ;
        RECT 141.815 176.965 145.035 176.980 ;
        RECT 141.365 176.515 145.035 176.965 ;
        RECT 125.145 174.065 125.545 174.115 ;
        RECT 110.195 173.815 140.795 174.065 ;
        RECT 125.145 173.065 125.545 173.115 ;
        RECT 110.195 172.815 140.795 173.065 ;
        RECT 109.965 168.015 110.195 172.610 ;
        RECT 120.255 168.015 120.485 172.610 ;
        RECT 130.545 168.015 130.775 172.610 ;
        RECT 139.395 171.365 139.795 171.665 ;
        RECT 139.495 168.715 139.695 171.365 ;
        RECT 139.395 168.415 139.795 168.715 ;
        RECT 140.835 168.015 141.065 172.610 ;
        RECT 141.365 171.765 141.625 176.515 ;
        RECT 141.815 176.500 145.035 176.515 ;
        RECT 143.855 176.165 144.300 176.170 ;
        RECT 142.495 176.090 142.895 176.115 ;
        RECT 142.485 175.790 142.930 176.090 ;
        RECT 143.845 175.870 144.300 176.165 ;
        RECT 143.845 175.865 144.295 175.870 ;
        RECT 142.075 175.315 142.520 175.365 ;
        RECT 142.045 175.065 142.520 175.315 ;
        RECT 143.445 175.065 143.900 175.365 ;
        RECT 142.045 174.465 142.495 175.065 ;
        RECT 142.045 174.415 142.445 174.465 ;
        RECT 141.815 174.165 144.575 174.260 ;
        RECT 141.815 173.815 144.595 174.165 ;
        RECT 141.815 173.780 144.575 173.815 ;
        RECT 143.595 172.915 143.995 173.215 ;
        RECT 142.595 171.915 143.045 172.265 ;
        RECT 143.695 172.175 143.845 172.915 ;
        RECT 143.625 171.945 143.915 172.175 ;
        RECT 141.365 171.740 142.045 171.765 ;
        RECT 141.365 171.320 142.205 171.740 ;
        RECT 142.455 171.725 142.685 171.740 ;
        RECT 142.935 171.725 143.165 171.740 ;
        RECT 142.385 171.325 142.685 171.725 ;
        RECT 142.925 171.325 143.225 171.725 ;
        RECT 142.455 171.320 142.685 171.325 ;
        RECT 142.935 171.320 143.165 171.325 ;
        RECT 143.415 171.320 143.645 171.740 ;
        RECT 143.895 171.565 144.125 171.740 ;
        RECT 143.895 171.415 144.645 171.565 ;
        RECT 143.895 171.320 144.125 171.415 ;
        RECT 141.365 171.315 142.045 171.320 ;
        RECT 141.365 170.665 141.625 171.315 ;
        RECT 142.095 170.815 142.495 171.115 ;
        RECT 141.295 170.365 141.695 170.665 ;
        RECT 141.365 169.665 141.625 170.365 ;
        RECT 142.195 170.095 142.445 170.815 ;
        RECT 143.145 170.165 143.445 171.115 ;
        RECT 144.495 170.665 144.645 171.415 ;
        RECT 144.845 171.365 145.245 171.665 ;
        RECT 144.395 170.365 144.795 170.665 ;
        RECT 142.185 169.865 142.475 170.095 ;
        RECT 143.095 169.865 143.495 170.165 ;
        RECT 141.365 169.660 142.045 169.665 ;
        RECT 141.365 169.240 142.205 169.660 ;
        RECT 142.385 169.265 142.685 169.665 ;
        RECT 142.925 169.265 143.225 169.665 ;
        RECT 142.455 169.240 142.685 169.265 ;
        RECT 142.935 169.240 143.165 169.265 ;
        RECT 143.415 169.240 143.645 169.660 ;
        RECT 143.895 169.515 144.125 169.660 ;
        RECT 144.495 169.515 144.645 170.365 ;
        RECT 143.895 169.365 144.645 169.515 ;
        RECT 143.895 169.240 144.125 169.365 ;
        RECT 141.365 169.215 142.045 169.240 ;
        RECT 141.365 168.815 141.625 169.215 ;
        RECT 141.365 168.015 141.645 168.815 ;
        RECT 142.595 168.715 143.045 169.065 ;
        RECT 143.625 168.805 143.915 169.035 ;
        RECT 143.695 168.115 143.845 168.805 ;
        RECT 77.465 161.340 77.765 161.590 ;
        RECT 83.015 161.590 107.790 161.740 ;
        RECT 109.245 166.315 141.645 168.015 ;
        RECT 143.545 167.815 143.945 168.115 ;
        RECT 141.945 167.195 142.395 167.715 ;
        RECT 144.395 167.365 144.795 167.665 ;
        RECT 141.935 166.835 142.395 167.195 ;
        RECT 143.645 166.865 144.045 167.165 ;
        RECT 141.945 166.815 142.395 166.835 ;
        RECT 142.695 166.365 143.095 166.665 ;
        RECT 143.745 166.525 143.895 166.865 ;
        RECT 109.245 161.865 109.745 166.315 ;
        RECT 109.965 162.610 110.195 166.315 ;
        RECT 120.255 162.610 120.485 166.315 ;
        RECT 130.545 162.610 130.775 166.315 ;
        RECT 140.835 162.610 141.065 166.315 ;
        RECT 142.725 166.295 143.015 166.365 ;
        RECT 143.685 166.295 143.975 166.525 ;
        RECT 142.440 165.735 142.745 166.135 ;
        RECT 142.980 165.735 143.280 166.135 ;
        RECT 142.515 165.715 142.745 165.735 ;
        RECT 142.995 165.715 143.225 165.735 ;
        RECT 143.475 165.715 143.705 166.135 ;
        RECT 143.955 166.015 144.185 166.135 ;
        RECT 144.445 166.015 144.645 167.365 ;
        RECT 143.955 165.865 144.645 166.015 ;
        RECT 143.955 165.715 144.185 165.865 ;
        RECT 143.195 165.115 143.495 165.565 ;
        RECT 143.145 164.815 143.545 165.115 ;
        RECT 143.195 164.315 143.495 164.815 ;
        RECT 143.205 164.305 143.495 164.315 ;
        RECT 142.515 164.135 142.745 164.145 ;
        RECT 142.995 164.135 143.225 164.145 ;
        RECT 142.440 163.735 142.745 164.135 ;
        RECT 142.980 163.735 143.280 164.135 ;
        RECT 142.515 163.725 142.745 163.735 ;
        RECT 142.995 163.725 143.225 163.735 ;
        RECT 143.475 163.725 143.705 164.145 ;
        RECT 143.955 164.015 144.185 164.145 ;
        RECT 144.445 164.015 144.645 165.865 ;
        RECT 144.945 166.065 145.095 171.365 ;
        RECT 145.445 170.215 145.595 179.965 ;
        RECT 145.895 175.365 146.045 180.515 ;
        RECT 145.795 175.065 146.195 175.365 ;
        RECT 145.845 173.265 146.145 173.665 ;
        RECT 145.895 172.265 146.045 173.265 ;
        RECT 145.795 171.965 146.195 172.265 ;
        RECT 145.245 169.915 145.645 170.215 ;
        RECT 145.245 169.315 145.645 169.615 ;
        RECT 144.945 165.765 145.345 166.065 ;
        RECT 145.495 164.115 145.645 169.315 ;
        RECT 145.895 169.015 146.045 171.965 ;
        RECT 145.795 168.715 146.195 169.015 ;
        RECT 146.345 168.115 146.495 183.165 ;
        RECT 146.695 182.715 147.095 183.015 ;
        RECT 146.745 173.165 146.895 182.715 ;
        RECT 147.095 181.450 147.495 181.750 ;
        RECT 147.195 174.715 147.345 181.450 ;
        RECT 147.645 177.915 147.795 184.490 ;
        RECT 148.090 181.240 148.240 184.490 ;
        RECT 147.940 180.940 148.340 181.240 ;
        RECT 148.895 179.615 149.245 185.065 ;
        RECT 150.165 184.390 150.315 184.415 ;
        RECT 150.040 184.090 150.440 184.390 ;
        RECT 148.845 179.265 149.295 179.615 ;
        RECT 147.995 178.715 148.395 179.015 ;
        RECT 147.545 177.515 147.845 177.915 ;
        RECT 147.095 174.415 147.495 174.715 ;
        RECT 146.645 172.865 147.045 173.165 ;
        RECT 146.145 167.815 146.545 168.115 ;
        RECT 145.795 166.465 146.195 166.765 ;
        RECT 143.955 163.865 144.645 164.015 ;
        RECT 143.955 163.725 144.185 163.865 ;
        RECT 145.345 163.815 145.745 164.115 ;
        RECT 145.895 163.565 146.045 166.465 ;
        RECT 142.725 163.515 143.015 163.565 ;
        RECT 142.645 163.215 143.045 163.515 ;
        RECT 143.685 163.335 143.975 163.565 ;
        RECT 143.745 162.865 143.895 163.335 ;
        RECT 145.795 163.265 146.195 163.565 ;
        RECT 146.345 162.865 146.495 167.815 ;
        RECT 146.745 167.215 146.895 172.865 ;
        RECT 146.645 166.915 147.045 167.215 ;
        RECT 147.195 165.065 147.345 174.415 ;
        RECT 147.645 171.215 147.795 177.515 ;
        RECT 148.095 173.615 148.245 178.715 ;
        RECT 148.445 178.115 148.745 178.515 ;
        RECT 147.945 173.315 148.345 173.615 ;
        RECT 148.495 171.715 148.645 178.115 ;
        RECT 148.895 174.165 149.245 179.265 ;
        RECT 148.845 173.815 149.295 174.165 ;
        RECT 148.395 171.665 148.645 171.715 ;
        RECT 148.245 171.365 148.645 171.665 ;
        RECT 147.545 170.815 147.845 171.215 ;
        RECT 148.495 166.715 148.645 171.365 ;
        RECT 148.895 167.115 149.245 173.815 ;
        RECT 148.295 166.415 148.695 166.715 ;
        RECT 147.095 164.765 147.495 165.065 ;
        RECT 143.595 162.565 143.995 162.865 ;
        RECT 146.095 162.565 146.495 162.865 ;
        RECT 110.195 162.115 140.895 162.415 ;
        RECT 83.015 161.340 83.315 161.590 ;
        RECT 109.245 161.515 141.445 161.865 ;
        RECT 105.190 161.190 105.590 161.240 ;
        RECT 150.215 161.190 150.365 184.090 ;
        RECT 105.190 161.040 150.365 161.190 ;
        RECT 105.190 160.940 105.590 161.040 ;
        RECT 30.165 160.465 142.115 160.615 ;
        RECT 20.205 159.800 37.535 160.185 ;
        RECT 20.205 159.705 26.600 159.800 ;
        RECT 10.815 159.215 11.415 159.365 ;
        RECT 10.240 158.540 10.640 158.840 ;
        RECT 10.815 155.765 10.965 159.215 ;
        RECT 20.220 158.805 20.585 159.110 ;
        RECT 20.355 158.640 20.585 158.805 ;
        RECT 20.220 158.440 20.585 158.640 ;
        RECT 23.245 158.870 23.550 158.920 ;
        RECT 23.715 158.870 24.020 158.920 ;
        RECT 24.210 158.875 24.655 159.705 ;
        RECT 24.795 158.875 25.025 159.160 ;
        RECT 23.245 158.640 24.065 158.870 ;
        RECT 23.245 158.560 23.550 158.640 ;
        RECT 23.715 158.560 24.020 158.640 ;
        RECT 20.220 158.335 20.580 158.440 ;
        RECT 20.205 156.985 23.885 157.465 ;
        RECT 23.505 155.980 23.735 156.050 ;
        RECT 21.580 155.825 21.885 155.880 ;
        RECT 22.050 155.825 22.355 155.880 ;
        RECT 21.580 155.765 22.400 155.825 ;
        RECT 10.815 155.615 22.400 155.765 ;
        RECT 23.465 155.675 23.825 155.980 ;
        RECT 21.580 155.595 22.400 155.615 ;
        RECT 21.580 155.520 21.885 155.595 ;
        RECT 22.050 155.520 22.355 155.595 ;
        RECT 23.505 155.510 23.735 155.675 ;
        RECT 24.210 155.610 25.025 158.875 ;
        RECT 25.275 157.010 25.505 159.160 ;
        RECT 25.755 158.845 25.985 159.160 ;
        RECT 26.290 158.845 26.600 159.705 ;
        RECT 28.395 159.705 37.535 159.800 ;
        RECT 27.095 159.300 27.400 159.660 ;
        RECT 27.565 159.300 27.870 159.660 ;
        RECT 25.230 156.705 25.590 157.010 ;
        RECT 25.275 156.540 25.505 156.705 ;
        RECT 25.230 156.235 25.590 156.540 ;
        RECT 23.465 155.205 23.825 155.510 ;
        RECT 21.585 154.460 23.885 154.745 ;
        RECT 24.210 154.460 24.655 155.610 ;
        RECT 24.795 155.160 25.025 155.610 ;
        RECT 25.275 155.160 25.505 156.235 ;
        RECT 25.755 155.610 26.600 158.845 ;
        RECT 26.895 158.225 27.125 159.160 ;
        RECT 26.810 157.920 27.170 158.225 ;
        RECT 26.895 157.755 27.125 157.920 ;
        RECT 26.810 157.450 27.170 157.755 ;
        RECT 25.755 155.160 25.985 155.610 ;
        RECT 24.985 154.660 25.760 155.020 ;
        RECT 26.290 154.460 26.600 155.610 ;
        RECT 26.895 155.160 27.125 157.450 ;
        RECT 27.375 156.960 27.605 159.160 ;
        RECT 27.855 158.225 28.085 159.160 ;
        RECT 28.395 158.810 28.715 159.705 ;
        RECT 28.995 158.810 29.225 159.160 ;
        RECT 27.800 157.920 28.160 158.225 ;
        RECT 27.855 157.755 28.085 157.920 ;
        RECT 27.800 157.450 28.160 157.755 ;
        RECT 27.280 156.655 27.640 156.960 ;
        RECT 27.375 156.490 27.605 156.655 ;
        RECT 27.280 156.185 27.640 156.490 ;
        RECT 27.375 155.160 27.605 156.185 ;
        RECT 27.855 155.160 28.085 157.450 ;
        RECT 28.395 155.380 29.225 158.810 ;
        RECT 29.475 156.140 29.705 159.160 ;
        RECT 29.955 158.800 30.185 159.160 ;
        RECT 30.515 158.800 31.305 159.705 ;
        RECT 31.975 159.140 32.835 159.370 ;
        RECT 29.430 155.835 29.790 156.140 ;
        RECT 29.475 155.670 29.705 155.835 ;
        RECT 28.395 154.460 28.715 155.380 ;
        RECT 28.995 155.160 29.225 155.380 ;
        RECT 29.430 155.365 29.790 155.670 ;
        RECT 29.955 155.380 31.305 158.800 ;
        RECT 31.695 158.760 31.925 158.980 ;
        RECT 31.630 158.455 31.990 158.760 ;
        RECT 31.695 158.290 31.925 158.455 ;
        RECT 31.630 157.985 31.990 158.290 ;
        RECT 29.475 155.160 29.705 155.365 ;
        RECT 29.955 155.160 30.185 155.380 ;
        RECT 29.170 154.660 29.945 155.020 ;
        RECT 30.515 154.460 31.305 155.380 ;
        RECT 31.695 154.980 31.925 157.985 ;
        RECT 32.885 157.770 33.115 158.980 ;
        RECT 32.820 157.465 33.180 157.770 ;
        RECT 32.885 157.300 33.115 157.465 ;
        RECT 32.820 156.995 33.180 157.300 ;
        RECT 32.885 154.980 33.115 156.995 ;
        RECT 21.585 154.100 31.305 154.460 ;
        RECT 31.635 154.310 33.230 154.820 ;
        RECT 33.435 154.100 33.875 159.705 ;
        RECT 34.505 159.140 35.365 159.370 ;
        RECT 35.695 159.140 36.555 159.370 ;
        RECT 34.225 157.780 34.455 158.980 ;
        RECT 34.160 157.475 34.520 157.780 ;
        RECT 34.225 157.310 34.455 157.475 ;
        RECT 34.160 157.005 34.520 157.310 ;
        RECT 34.225 154.980 34.455 157.005 ;
        RECT 35.415 156.140 35.645 158.980 ;
        RECT 36.605 157.780 36.835 158.980 ;
        RECT 36.540 157.475 36.900 157.780 ;
        RECT 36.605 157.310 36.835 157.475 ;
        RECT 36.540 157.005 36.900 157.310 ;
        RECT 35.350 155.835 35.710 156.140 ;
        RECT 35.415 155.670 35.645 155.835 ;
        RECT 35.350 155.365 35.710 155.670 ;
        RECT 35.415 154.980 35.645 155.365 ;
        RECT 36.605 154.980 36.835 157.005 ;
        RECT 34.505 154.790 35.365 154.820 ;
        RECT 35.695 154.790 36.555 154.820 ;
        RECT 34.505 154.310 36.555 154.790 ;
        RECT 37.145 154.100 37.535 159.705 ;
        RECT 21.585 153.690 37.535 154.100 ;
        RECT 37.715 159.795 74.610 160.190 ;
        RECT 37.715 159.705 41.175 159.795 ;
        RECT 37.715 154.505 38.200 159.705 ;
        RECT 38.435 158.650 38.665 159.115 ;
        RECT 38.370 158.345 38.730 158.650 ;
        RECT 38.435 158.180 38.665 158.345 ;
        RECT 38.370 157.875 38.730 158.180 ;
        RECT 38.435 155.115 38.665 157.875 ;
        RECT 38.915 157.620 39.145 159.115 ;
        RECT 39.395 158.650 39.625 159.115 ;
        RECT 39.330 158.345 39.690 158.650 ;
        RECT 39.395 158.180 39.625 158.345 ;
        RECT 39.330 157.875 39.690 158.180 ;
        RECT 38.810 157.315 39.170 157.620 ;
        RECT 38.915 157.150 39.145 157.315 ;
        RECT 38.810 156.845 39.170 157.150 ;
        RECT 38.915 155.115 39.145 156.845 ;
        RECT 39.395 155.115 39.625 157.875 ;
        RECT 39.875 157.620 40.105 159.115 ;
        RECT 40.355 158.650 40.585 159.115 ;
        RECT 40.820 158.650 41.175 159.705 ;
        RECT 42.395 159.705 74.610 159.795 ;
        RECT 41.445 159.550 41.750 159.615 ;
        RECT 41.915 159.550 42.220 159.615 ;
        RECT 41.445 159.320 42.220 159.550 ;
        RECT 41.445 159.255 41.750 159.320 ;
        RECT 41.915 159.255 42.220 159.320 ;
        RECT 41.495 158.880 41.725 159.115 ;
        RECT 40.290 158.345 41.175 158.650 ;
        RECT 40.315 158.180 41.175 158.345 ;
        RECT 40.290 157.875 41.175 158.180 ;
        RECT 40.315 157.870 41.175 157.875 ;
        RECT 39.770 157.315 40.130 157.620 ;
        RECT 39.875 157.150 40.105 157.315 ;
        RECT 39.770 156.845 40.130 157.150 ;
        RECT 39.875 155.115 40.105 156.845 ;
        RECT 40.355 155.115 40.585 157.870 ;
        RECT 40.820 157.830 41.175 157.870 ;
        RECT 41.385 158.115 41.725 158.880 ;
        RECT 41.935 159.000 42.165 159.115 ;
        RECT 42.395 159.000 42.880 159.705 ;
        RECT 43.955 159.550 44.260 159.560 ;
        RECT 44.425 159.550 44.730 159.560 ;
        RECT 43.355 159.320 73.610 159.550 ;
        RECT 43.955 159.200 44.260 159.320 ;
        RECT 44.425 159.200 44.730 159.320 ;
        RECT 55.335 159.190 55.640 159.320 ;
        RECT 55.805 159.190 56.110 159.320 ;
        RECT 61.235 159.190 61.540 159.320 ;
        RECT 61.705 159.190 62.010 159.320 ;
        RECT 70.095 159.190 70.400 159.320 ;
        RECT 70.565 159.190 70.870 159.320 ;
        RECT 41.935 158.455 42.880 159.000 ;
        RECT 43.075 158.455 43.305 159.115 ;
        RECT 58.365 158.455 58.595 159.115 ;
        RECT 73.655 158.455 73.885 159.115 ;
        RECT 74.125 158.455 74.610 159.705 ;
        RECT 41.935 158.260 74.610 158.455 ;
        RECT 41.935 158.115 42.165 158.260 ;
        RECT 38.910 154.910 39.215 154.975 ;
        RECT 39.380 154.910 39.685 154.975 ;
        RECT 40.820 154.930 41.185 157.830 ;
        RECT 41.385 155.910 41.635 158.115 ;
        RECT 42.395 157.370 74.610 158.260 ;
        RECT 42.385 156.310 74.610 157.370 ;
        RECT 41.330 155.605 41.690 155.910 ;
        RECT 41.385 155.440 41.635 155.605 ;
        RECT 41.330 155.135 41.690 155.440 ;
        RECT 42.385 154.930 42.880 156.310 ;
        RECT 43.075 155.365 43.305 156.310 ;
        RECT 58.365 155.365 58.595 156.310 ;
        RECT 73.655 155.365 73.885 156.310 ;
        RECT 43.935 155.160 44.240 155.290 ;
        RECT 44.405 155.160 44.710 155.290 ;
        RECT 55.285 155.160 55.590 155.290 ;
        RECT 55.755 155.160 56.060 155.290 ;
        RECT 61.185 155.160 61.490 155.290 ;
        RECT 61.655 155.160 61.960 155.290 ;
        RECT 70.085 155.160 70.390 155.290 ;
        RECT 70.555 155.160 70.860 155.290 ;
        RECT 43.355 154.930 73.610 155.160 ;
        RECT 38.645 154.680 39.895 154.910 ;
        RECT 38.910 154.615 39.215 154.680 ;
        RECT 39.380 154.615 39.685 154.680 ;
        RECT 40.820 154.505 42.880 154.930 ;
        RECT 43.365 154.620 58.170 154.930 ;
        RECT 58.710 154.620 73.515 154.930 ;
        RECT 37.715 154.300 38.485 154.505 ;
        RECT 40.050 154.300 42.880 154.505 ;
        RECT 43.355 154.390 58.315 154.620 ;
        RECT 58.645 154.390 73.605 154.620 ;
        RECT 37.715 154.020 42.880 154.300 ;
        RECT 9.915 153.190 10.215 153.590 ;
        RECT 42.385 153.435 42.880 154.020 ;
        RECT 43.075 153.435 43.305 154.185 ;
        RECT 58.365 153.435 58.595 154.185 ;
        RECT 73.655 153.435 73.885 154.185 ;
        RECT 74.125 153.435 74.610 156.310 ;
        RECT 18.565 153.015 18.865 153.140 ;
        RECT 9.615 152.865 18.865 153.015 ;
        RECT 18.565 152.740 18.865 152.865 ;
        RECT 23.590 152.565 23.990 152.640 ;
        RECT 9.315 152.415 23.990 152.565 ;
        RECT 23.590 152.340 23.990 152.415 ;
        RECT 26.190 152.115 26.590 152.190 ;
        RECT 9.015 151.965 26.590 152.115 ;
        RECT 26.190 151.890 26.590 151.965 ;
        RECT 27.440 151.665 27.840 151.740 ;
        RECT 8.715 151.515 27.840 151.665 ;
        RECT 27.440 151.440 27.840 151.515 ;
        RECT 42.385 151.290 74.610 153.435 ;
        RECT 28.640 151.215 29.040 151.290 ;
        RECT 8.415 151.065 29.040 151.215 ;
        RECT 28.640 150.990 29.040 151.065 ;
        RECT 29.890 150.765 30.290 150.840 ;
        RECT 8.115 150.615 30.290 150.765 ;
        RECT 29.890 150.540 30.290 150.615 ;
        RECT 31.090 150.315 31.490 150.390 ;
        RECT 7.815 150.165 31.490 150.315 ;
        RECT 31.090 150.090 31.490 150.165 ;
        RECT 32.290 149.865 32.690 149.940 ;
        RECT 7.515 149.715 32.690 149.865 ;
        RECT 32.290 149.640 32.690 149.715 ;
        RECT 42.385 149.845 42.880 151.290 ;
        RECT 43.075 150.435 43.305 151.290 ;
        RECT 58.365 150.435 58.595 151.290 ;
        RECT 73.655 150.435 73.885 151.290 ;
        RECT 43.835 150.230 44.735 150.330 ;
        RECT 55.235 150.230 56.085 150.380 ;
        RECT 61.135 150.230 61.985 150.380 ;
        RECT 70.085 150.230 70.935 150.380 ;
        RECT 43.355 150.000 58.315 150.230 ;
        RECT 58.645 150.000 73.605 150.230 ;
        RECT 74.125 149.845 74.610 151.290 ;
        RECT 33.540 149.415 33.940 149.490 ;
        RECT 7.215 149.265 33.940 149.415 ;
        RECT 42.385 149.360 74.610 149.845 ;
        RECT 86.505 159.795 123.400 160.190 ;
        RECT 86.505 159.705 118.720 159.795 ;
        RECT 86.505 158.455 86.990 159.705 ;
        RECT 116.385 159.550 116.690 159.560 ;
        RECT 116.855 159.550 117.160 159.560 ;
        RECT 87.505 159.320 117.760 159.550 ;
        RECT 90.245 159.190 90.550 159.320 ;
        RECT 90.715 159.190 91.020 159.320 ;
        RECT 99.105 159.190 99.410 159.320 ;
        RECT 99.575 159.190 99.880 159.320 ;
        RECT 105.005 159.190 105.310 159.320 ;
        RECT 105.475 159.190 105.780 159.320 ;
        RECT 116.385 159.200 116.690 159.320 ;
        RECT 116.855 159.200 117.160 159.320 ;
        RECT 87.230 158.455 87.460 159.115 ;
        RECT 102.520 158.455 102.750 159.115 ;
        RECT 117.810 158.455 118.040 159.115 ;
        RECT 118.235 159.000 118.720 159.705 ;
        RECT 119.940 159.705 123.400 159.795 ;
        RECT 118.895 159.550 119.200 159.615 ;
        RECT 119.365 159.550 119.670 159.615 ;
        RECT 118.895 159.320 119.670 159.550 ;
        RECT 118.895 159.255 119.200 159.320 ;
        RECT 119.365 159.255 119.670 159.320 ;
        RECT 118.950 159.000 119.180 159.115 ;
        RECT 118.235 158.455 119.180 159.000 ;
        RECT 86.505 158.260 119.180 158.455 ;
        RECT 86.505 157.370 118.720 158.260 ;
        RECT 118.950 158.115 119.180 158.260 ;
        RECT 119.390 158.880 119.620 159.115 ;
        RECT 119.390 158.115 119.730 158.880 ;
        RECT 86.505 156.310 118.730 157.370 ;
        RECT 86.505 153.435 86.990 156.310 ;
        RECT 87.230 155.365 87.460 156.310 ;
        RECT 102.520 155.365 102.750 156.310 ;
        RECT 117.810 155.365 118.040 156.310 ;
        RECT 90.255 155.160 90.560 155.290 ;
        RECT 90.725 155.160 91.030 155.290 ;
        RECT 99.155 155.160 99.460 155.290 ;
        RECT 99.625 155.160 99.930 155.290 ;
        RECT 105.055 155.160 105.360 155.290 ;
        RECT 105.525 155.160 105.830 155.290 ;
        RECT 116.405 155.160 116.710 155.290 ;
        RECT 116.875 155.160 117.180 155.290 ;
        RECT 87.505 154.930 117.760 155.160 ;
        RECT 118.235 154.930 118.730 156.310 ;
        RECT 119.480 155.910 119.730 158.115 ;
        RECT 119.940 158.650 120.295 159.705 ;
        RECT 120.530 158.650 120.760 159.115 ;
        RECT 119.940 158.345 120.825 158.650 ;
        RECT 119.940 158.180 120.800 158.345 ;
        RECT 119.940 157.875 120.825 158.180 ;
        RECT 119.940 157.870 120.800 157.875 ;
        RECT 119.940 157.830 120.295 157.870 ;
        RECT 119.425 155.605 119.785 155.910 ;
        RECT 119.480 155.440 119.730 155.605 ;
        RECT 119.425 155.135 119.785 155.440 ;
        RECT 119.930 154.930 120.295 157.830 ;
        RECT 120.530 155.115 120.760 157.870 ;
        RECT 121.010 157.620 121.240 159.115 ;
        RECT 121.490 158.650 121.720 159.115 ;
        RECT 121.425 158.345 121.785 158.650 ;
        RECT 121.490 158.180 121.720 158.345 ;
        RECT 121.425 157.875 121.785 158.180 ;
        RECT 120.985 157.315 121.345 157.620 ;
        RECT 121.010 157.150 121.240 157.315 ;
        RECT 120.985 156.845 121.345 157.150 ;
        RECT 121.010 155.115 121.240 156.845 ;
        RECT 121.490 155.115 121.720 157.875 ;
        RECT 121.970 157.620 122.200 159.115 ;
        RECT 122.450 158.650 122.680 159.115 ;
        RECT 122.385 158.345 122.745 158.650 ;
        RECT 122.450 158.180 122.680 158.345 ;
        RECT 122.385 157.875 122.745 158.180 ;
        RECT 121.945 157.315 122.305 157.620 ;
        RECT 121.970 157.150 122.200 157.315 ;
        RECT 121.945 156.845 122.305 157.150 ;
        RECT 121.970 155.115 122.200 156.845 ;
        RECT 122.450 155.115 122.680 157.875 ;
        RECT 87.600 154.620 102.405 154.930 ;
        RECT 102.945 154.620 117.750 154.930 ;
        RECT 87.510 154.390 102.470 154.620 ;
        RECT 102.800 154.390 117.760 154.620 ;
        RECT 118.235 154.505 120.295 154.930 ;
        RECT 121.430 154.910 121.735 154.975 ;
        RECT 121.900 154.910 122.205 154.975 ;
        RECT 121.220 154.680 122.470 154.910 ;
        RECT 121.430 154.615 121.735 154.680 ;
        RECT 121.900 154.615 122.205 154.680 ;
        RECT 122.915 154.505 123.400 159.705 ;
        RECT 118.235 154.300 121.065 154.505 ;
        RECT 122.630 154.300 123.400 154.505 ;
        RECT 87.230 153.435 87.460 154.185 ;
        RECT 102.520 153.435 102.750 154.185 ;
        RECT 117.810 153.435 118.040 154.185 ;
        RECT 118.235 154.020 123.400 154.300 ;
        RECT 123.580 159.800 140.910 160.185 ;
        RECT 123.580 159.705 132.720 159.800 ;
        RECT 123.580 154.100 123.970 159.705 ;
        RECT 124.560 159.140 125.420 159.370 ;
        RECT 125.750 159.140 126.610 159.370 ;
        RECT 124.280 157.780 124.510 158.980 ;
        RECT 124.215 157.475 124.575 157.780 ;
        RECT 124.280 157.310 124.510 157.475 ;
        RECT 124.215 157.005 124.575 157.310 ;
        RECT 124.280 154.980 124.510 157.005 ;
        RECT 125.470 156.140 125.700 158.980 ;
        RECT 126.660 157.780 126.890 158.980 ;
        RECT 126.595 157.475 126.955 157.780 ;
        RECT 126.660 157.310 126.890 157.475 ;
        RECT 126.595 157.005 126.955 157.310 ;
        RECT 125.405 155.835 125.765 156.140 ;
        RECT 125.470 155.670 125.700 155.835 ;
        RECT 125.405 155.365 125.765 155.670 ;
        RECT 125.470 154.980 125.700 155.365 ;
        RECT 126.660 154.980 126.890 157.005 ;
        RECT 124.560 154.790 125.420 154.820 ;
        RECT 125.750 154.790 126.610 154.820 ;
        RECT 124.560 154.310 126.610 154.790 ;
        RECT 127.240 154.100 127.680 159.705 ;
        RECT 128.280 159.140 129.140 159.370 ;
        RECT 128.000 157.770 128.230 158.980 ;
        RECT 129.190 158.760 129.420 158.980 ;
        RECT 129.810 158.800 130.600 159.705 ;
        RECT 130.930 158.800 131.160 159.160 ;
        RECT 129.125 158.455 129.485 158.760 ;
        RECT 129.190 158.290 129.420 158.455 ;
        RECT 129.125 157.985 129.485 158.290 ;
        RECT 127.935 157.465 128.295 157.770 ;
        RECT 128.000 157.300 128.230 157.465 ;
        RECT 127.935 156.995 128.295 157.300 ;
        RECT 128.000 154.980 128.230 156.995 ;
        RECT 129.190 154.980 129.420 157.985 ;
        RECT 129.810 155.380 131.160 158.800 ;
        RECT 131.410 156.140 131.640 159.160 ;
        RECT 131.890 158.810 132.120 159.160 ;
        RECT 132.400 158.810 132.720 159.705 ;
        RECT 134.515 159.705 140.910 159.800 ;
        RECT 133.245 159.300 133.550 159.660 ;
        RECT 133.715 159.300 134.020 159.660 ;
        RECT 131.325 155.835 131.685 156.140 ;
        RECT 131.410 155.670 131.640 155.835 ;
        RECT 127.885 154.310 129.480 154.820 ;
        RECT 129.810 154.460 130.600 155.380 ;
        RECT 130.930 155.160 131.160 155.380 ;
        RECT 131.325 155.365 131.685 155.670 ;
        RECT 131.890 155.380 132.720 158.810 ;
        RECT 133.030 158.225 133.260 159.160 ;
        RECT 132.955 157.920 133.315 158.225 ;
        RECT 133.030 157.755 133.260 157.920 ;
        RECT 132.955 157.450 133.315 157.755 ;
        RECT 131.410 155.160 131.640 155.365 ;
        RECT 131.890 155.160 132.120 155.380 ;
        RECT 131.170 154.660 131.945 155.020 ;
        RECT 132.400 154.460 132.720 155.380 ;
        RECT 133.030 155.160 133.260 157.450 ;
        RECT 133.510 156.960 133.740 159.160 ;
        RECT 133.990 158.225 134.220 159.160 ;
        RECT 134.515 158.845 134.825 159.705 ;
        RECT 135.130 158.845 135.360 159.160 ;
        RECT 133.945 157.920 134.305 158.225 ;
        RECT 133.990 157.755 134.220 157.920 ;
        RECT 133.945 157.450 134.305 157.755 ;
        RECT 133.475 156.655 133.835 156.960 ;
        RECT 133.510 156.490 133.740 156.655 ;
        RECT 133.475 156.185 133.835 156.490 ;
        RECT 133.510 155.160 133.740 156.185 ;
        RECT 133.990 155.160 134.220 157.450 ;
        RECT 134.515 155.610 135.360 158.845 ;
        RECT 135.610 157.010 135.840 159.160 ;
        RECT 136.090 158.875 136.320 159.160 ;
        RECT 136.460 158.875 136.905 159.705 ;
        RECT 135.525 156.705 135.885 157.010 ;
        RECT 135.610 156.540 135.840 156.705 ;
        RECT 135.525 156.235 135.885 156.540 ;
        RECT 134.515 154.460 134.825 155.610 ;
        RECT 135.130 155.160 135.360 155.610 ;
        RECT 135.610 155.160 135.840 156.235 ;
        RECT 136.090 155.610 136.905 158.875 ;
        RECT 137.095 158.870 137.400 158.920 ;
        RECT 137.565 158.870 137.870 158.920 ;
        RECT 137.050 158.640 137.870 158.870 ;
        RECT 137.095 158.560 137.400 158.640 ;
        RECT 137.565 158.560 137.870 158.640 ;
        RECT 140.530 158.805 140.895 159.110 ;
        RECT 140.530 158.640 140.760 158.805 ;
        RECT 140.530 158.440 140.895 158.640 ;
        RECT 140.535 158.335 140.895 158.440 ;
        RECT 137.230 156.985 140.910 157.465 ;
        RECT 137.380 155.980 137.610 156.050 ;
        RECT 137.290 155.675 137.650 155.980 ;
        RECT 138.760 155.825 139.065 155.880 ;
        RECT 139.230 155.825 139.535 155.880 ;
        RECT 138.715 155.765 139.535 155.825 ;
        RECT 141.965 155.765 142.115 160.465 ;
        RECT 150.600 158.840 150.750 219.290 ;
        RECT 151.000 217.990 151.300 218.390 ;
        RECT 150.475 158.540 150.875 158.840 ;
        RECT 136.090 155.160 136.320 155.610 ;
        RECT 135.355 154.660 136.130 155.020 ;
        RECT 136.460 154.460 136.905 155.610 ;
        RECT 137.380 155.510 137.610 155.675 ;
        RECT 138.715 155.615 142.115 155.765 ;
        RECT 138.715 155.595 139.535 155.615 ;
        RECT 138.760 155.520 139.065 155.595 ;
        RECT 139.230 155.520 139.535 155.595 ;
        RECT 137.290 155.205 137.650 155.510 ;
        RECT 137.230 154.460 139.530 154.745 ;
        RECT 129.810 154.100 139.530 154.460 ;
        RECT 118.235 153.435 118.730 154.020 ;
        RECT 123.580 153.690 139.530 154.100 ;
        RECT 151.050 153.590 151.200 217.990 ;
        RECT 86.505 151.290 118.730 153.435 ;
        RECT 150.900 153.190 151.200 153.590 ;
        RECT 151.350 216.640 151.650 217.040 ;
        RECT 142.250 153.015 142.550 153.140 ;
        RECT 151.350 153.015 151.500 216.640 ;
        RECT 142.250 152.865 151.500 153.015 ;
        RECT 151.650 215.240 151.950 215.640 ;
        RECT 142.250 152.740 142.550 152.865 ;
        RECT 137.125 152.565 137.525 152.640 ;
        RECT 151.650 152.565 151.800 215.240 ;
        RECT 137.125 152.415 151.800 152.565 ;
        RECT 151.950 213.890 152.250 214.290 ;
        RECT 137.125 152.340 137.525 152.415 ;
        RECT 134.525 152.115 134.925 152.190 ;
        RECT 151.950 152.115 152.100 213.890 ;
        RECT 134.525 151.965 152.100 152.115 ;
        RECT 152.250 212.490 152.550 212.890 ;
        RECT 134.525 151.890 134.925 151.965 ;
        RECT 133.275 151.665 133.675 151.740 ;
        RECT 152.250 151.665 152.400 212.490 ;
        RECT 133.275 151.515 152.400 151.665 ;
        RECT 152.550 211.190 152.850 211.590 ;
        RECT 133.275 151.440 133.675 151.515 ;
        RECT 86.505 149.845 86.990 151.290 ;
        RECT 87.230 150.435 87.460 151.290 ;
        RECT 102.520 150.435 102.750 151.290 ;
        RECT 117.810 150.435 118.040 151.290 ;
        RECT 90.180 150.230 91.030 150.380 ;
        RECT 99.130 150.230 99.980 150.380 ;
        RECT 105.030 150.230 105.880 150.380 ;
        RECT 116.380 150.230 117.280 150.330 ;
        RECT 87.510 150.000 102.470 150.230 ;
        RECT 102.800 150.000 117.760 150.230 ;
        RECT 118.235 149.845 118.730 151.290 ;
        RECT 132.075 151.215 132.475 151.290 ;
        RECT 152.550 151.215 152.700 211.190 ;
        RECT 132.075 151.065 152.700 151.215 ;
        RECT 152.850 209.840 153.150 210.240 ;
        RECT 132.075 150.990 132.475 151.065 ;
        RECT 130.825 150.765 131.225 150.840 ;
        RECT 152.850 150.765 153.000 209.840 ;
        RECT 130.825 150.615 153.000 150.765 ;
        RECT 153.150 208.440 153.450 208.840 ;
        RECT 130.825 150.540 131.225 150.615 ;
        RECT 129.625 150.315 130.025 150.390 ;
        RECT 153.150 150.315 153.300 208.440 ;
        RECT 129.625 150.165 153.300 150.315 ;
        RECT 153.450 207.090 153.750 207.490 ;
        RECT 129.625 150.090 130.025 150.165 ;
        RECT 86.505 149.360 118.730 149.845 ;
        RECT 128.425 149.865 128.825 149.940 ;
        RECT 153.450 149.865 153.600 207.090 ;
        RECT 128.425 149.715 153.600 149.865 ;
        RECT 153.750 205.790 154.050 206.190 ;
        RECT 128.425 149.640 128.825 149.715 ;
        RECT 127.175 149.415 127.575 149.490 ;
        RECT 153.750 149.415 153.900 205.790 ;
        RECT 33.540 149.190 33.940 149.265 ;
        RECT 127.175 149.265 153.900 149.415 ;
        RECT 154.050 204.390 154.350 204.790 ;
        RECT 127.175 149.190 127.575 149.265 ;
        RECT 34.690 148.965 35.090 149.040 ;
        RECT 6.915 148.815 35.090 148.965 ;
        RECT 34.690 148.740 35.090 148.815 ;
        RECT 47.290 148.965 47.690 149.040 ;
        RECT 82.890 148.965 83.290 149.040 ;
        RECT 113.425 148.965 113.825 149.040 ;
        RECT 47.290 148.815 113.825 148.965 ;
        RECT 47.290 148.740 47.690 148.815 ;
        RECT 82.890 148.740 83.290 148.815 ;
        RECT 113.425 148.740 113.825 148.815 ;
        RECT 126.025 148.965 126.425 149.040 ;
        RECT 154.050 148.965 154.200 204.390 ;
        RECT 126.025 148.815 154.200 148.965 ;
        RECT 154.350 203.040 154.650 203.440 ;
        RECT 126.025 148.740 126.425 148.815 ;
        RECT 37.440 148.515 37.840 148.590 ;
        RECT 6.615 148.365 37.840 148.515 ;
        RECT 37.440 148.290 37.840 148.365 ;
        RECT 51.140 148.515 51.540 148.590 ;
        RECT 82.440 148.515 82.840 148.590 ;
        RECT 109.575 148.515 109.975 148.590 ;
        RECT 51.140 148.365 109.975 148.515 ;
        RECT 51.140 148.290 51.540 148.365 ;
        RECT 82.440 148.290 82.840 148.365 ;
        RECT 109.575 148.290 109.975 148.365 ;
        RECT 123.275 148.515 123.675 148.590 ;
        RECT 154.350 148.515 154.500 203.040 ;
        RECT 123.275 148.365 154.500 148.515 ;
        RECT 154.650 201.640 154.950 202.040 ;
        RECT 123.275 148.290 123.675 148.365 ;
        RECT 41.290 148.065 41.690 148.140 ;
        RECT 6.315 147.915 41.690 148.065 ;
        RECT 41.290 147.840 41.690 147.915 ;
        RECT 54.990 148.065 55.390 148.140 ;
        RECT 81.990 148.065 82.390 148.140 ;
        RECT 105.725 148.065 106.125 148.140 ;
        RECT 54.990 147.915 106.125 148.065 ;
        RECT 54.990 147.840 55.390 147.915 ;
        RECT 81.990 147.840 82.390 147.915 ;
        RECT 105.725 147.840 106.125 147.915 ;
        RECT 119.425 148.065 119.825 148.140 ;
        RECT 154.650 148.065 154.800 201.640 ;
        RECT 119.425 147.915 154.800 148.065 ;
        RECT 154.950 200.340 155.250 200.740 ;
        RECT 119.425 147.840 119.825 147.915 ;
        RECT 43.240 147.615 43.640 147.690 ;
        RECT 6.015 147.465 43.640 147.615 ;
        RECT 43.240 147.390 43.640 147.465 ;
        RECT 56.890 147.615 57.290 147.690 ;
        RECT 81.540 147.615 81.940 147.690 ;
        RECT 103.825 147.615 104.225 147.690 ;
        RECT 56.890 147.465 104.225 147.615 ;
        RECT 56.890 147.390 57.290 147.465 ;
        RECT 81.540 147.390 81.940 147.465 ;
        RECT 103.825 147.390 104.225 147.465 ;
        RECT 117.475 147.615 117.875 147.690 ;
        RECT 154.950 147.615 155.100 200.340 ;
        RECT 117.475 147.465 155.100 147.615 ;
        RECT 155.250 198.990 155.550 199.390 ;
        RECT 117.475 147.390 117.875 147.465 ;
        RECT 44.090 147.165 44.490 147.240 ;
        RECT 5.715 147.015 44.490 147.165 ;
        RECT 44.090 146.940 44.490 147.015 ;
        RECT 57.840 147.165 58.240 147.240 ;
        RECT 81.090 147.165 81.490 147.240 ;
        RECT 102.875 147.165 103.275 147.240 ;
        RECT 57.840 147.015 103.275 147.165 ;
        RECT 57.840 146.940 58.240 147.015 ;
        RECT 81.090 146.940 81.490 147.015 ;
        RECT 102.875 146.940 103.275 147.015 ;
        RECT 116.625 147.165 117.025 147.240 ;
        RECT 155.250 147.165 155.400 198.990 ;
        RECT 116.625 147.015 155.400 147.165 ;
        RECT 155.550 197.640 155.850 198.040 ;
        RECT 116.625 146.940 117.025 147.015 ;
        RECT 36.540 146.715 36.940 146.790 ;
        RECT 45.190 146.715 45.590 146.790 ;
        RECT 36.540 146.565 45.590 146.715 ;
        RECT 36.540 146.490 36.940 146.565 ;
        RECT 45.190 146.490 45.590 146.565 ;
        RECT 65.290 146.715 65.690 146.790 ;
        RECT 80.640 146.715 81.040 146.790 ;
        RECT 95.425 146.715 95.825 146.790 ;
        RECT 65.290 146.565 95.825 146.715 ;
        RECT 65.290 146.490 65.690 146.565 ;
        RECT 80.640 146.490 81.040 146.565 ;
        RECT 95.425 146.490 95.825 146.565 ;
        RECT 115.525 146.715 115.925 146.790 ;
        RECT 124.175 146.715 124.575 146.790 ;
        RECT 115.525 146.565 124.575 146.715 ;
        RECT 115.525 146.490 115.925 146.565 ;
        RECT 124.175 146.490 124.575 146.565 ;
        RECT 58.890 146.265 59.290 146.340 ;
        RECT 5.415 146.115 59.290 146.265 ;
        RECT 58.890 146.040 59.290 146.115 ;
        RECT 66.090 146.265 66.490 146.340 ;
        RECT 80.190 146.265 80.590 146.340 ;
        RECT 94.625 146.265 95.025 146.340 ;
        RECT 66.090 146.115 95.025 146.265 ;
        RECT 66.090 146.040 66.490 146.115 ;
        RECT 80.190 146.040 80.590 146.115 ;
        RECT 94.625 146.040 95.025 146.115 ;
        RECT 101.825 146.265 102.225 146.340 ;
        RECT 155.550 146.265 155.700 197.640 ;
        RECT 101.825 146.115 155.700 146.265 ;
        RECT 155.850 196.190 156.150 196.590 ;
        RECT 101.825 146.040 102.225 146.115 ;
        RECT 59.840 145.815 60.240 145.890 ;
        RECT 5.115 145.665 60.240 145.815 ;
        RECT 59.840 145.590 60.240 145.665 ;
        RECT 66.890 145.815 67.290 145.890 ;
        RECT 79.740 145.815 80.140 145.890 ;
        RECT 93.825 145.815 94.225 145.890 ;
        RECT 66.890 145.665 94.225 145.815 ;
        RECT 66.890 145.590 67.290 145.665 ;
        RECT 79.740 145.590 80.140 145.665 ;
        RECT 93.825 145.590 94.225 145.665 ;
        RECT 100.875 145.815 101.275 145.890 ;
        RECT 155.850 145.815 156.000 196.190 ;
        RECT 100.875 145.665 156.000 145.815 ;
        RECT 156.150 194.840 156.450 195.240 ;
        RECT 100.875 145.590 101.275 145.665 ;
        RECT 60.440 145.365 60.840 145.440 ;
        RECT 4.815 145.215 60.840 145.365 ;
        RECT 60.440 145.140 60.840 145.215 ;
        RECT 67.690 145.365 68.090 145.440 ;
        RECT 79.290 145.365 79.690 145.440 ;
        RECT 93.025 145.365 93.425 145.440 ;
        RECT 67.690 145.215 93.425 145.365 ;
        RECT 67.690 145.140 68.090 145.215 ;
        RECT 79.290 145.140 79.690 145.215 ;
        RECT 93.025 145.140 93.425 145.215 ;
        RECT 100.275 145.365 100.675 145.440 ;
        RECT 156.150 145.365 156.300 194.840 ;
        RECT 100.275 145.215 156.300 145.365 ;
        RECT 156.450 193.540 156.750 193.940 ;
        RECT 100.275 145.140 100.675 145.215 ;
        RECT 61.490 144.915 61.890 144.990 ;
        RECT 4.515 144.765 61.890 144.915 ;
        RECT 61.490 144.690 61.890 144.765 ;
        RECT 65.690 144.915 66.090 144.990 ;
        RECT 78.840 144.915 79.240 144.990 ;
        RECT 95.025 144.915 95.425 144.990 ;
        RECT 65.690 144.765 95.425 144.915 ;
        RECT 65.690 144.690 66.090 144.765 ;
        RECT 78.840 144.690 79.240 144.765 ;
        RECT 95.025 144.690 95.425 144.765 ;
        RECT 99.225 144.915 99.625 144.990 ;
        RECT 156.450 144.915 156.600 193.540 ;
        RECT 99.225 144.765 156.600 144.915 ;
        RECT 156.750 192.090 157.050 192.490 ;
        RECT 99.225 144.690 99.625 144.765 ;
        RECT 62.540 144.465 62.940 144.540 ;
        RECT 4.215 144.315 62.940 144.465 ;
        RECT 62.540 144.240 62.940 144.315 ;
        RECT 66.490 144.465 66.890 144.540 ;
        RECT 78.390 144.465 78.790 144.540 ;
        RECT 94.225 144.465 94.625 144.540 ;
        RECT 66.490 144.315 94.625 144.465 ;
        RECT 66.490 144.240 66.890 144.315 ;
        RECT 78.390 144.240 78.790 144.315 ;
        RECT 94.225 144.240 94.625 144.315 ;
        RECT 98.175 144.465 98.575 144.540 ;
        RECT 156.750 144.465 156.900 192.090 ;
        RECT 98.175 144.315 156.900 144.465 ;
        RECT 157.050 190.740 157.350 191.140 ;
        RECT 98.175 144.240 98.575 144.315 ;
        RECT 63.590 144.015 63.990 144.090 ;
        RECT 3.915 143.865 63.990 144.015 ;
        RECT 63.590 143.790 63.990 143.865 ;
        RECT 67.290 144.015 67.690 144.090 ;
        RECT 77.940 144.015 78.340 144.090 ;
        RECT 93.425 144.015 93.825 144.090 ;
        RECT 67.290 143.865 93.825 144.015 ;
        RECT 67.290 143.790 67.690 143.865 ;
        RECT 77.940 143.790 78.340 143.865 ;
        RECT 93.425 143.790 93.825 143.865 ;
        RECT 97.125 144.015 97.525 144.090 ;
        RECT 157.050 144.015 157.200 190.740 ;
        RECT 97.125 143.865 157.200 144.015 ;
        RECT 157.350 189.340 157.650 189.740 ;
        RECT 97.125 143.790 97.525 143.865 ;
        RECT 64.640 143.565 65.040 143.640 ;
        RECT 3.615 143.415 65.040 143.565 ;
        RECT 64.640 143.340 65.040 143.415 ;
        RECT 68.090 143.565 68.490 143.640 ;
        RECT 77.490 143.565 77.890 143.640 ;
        RECT 92.625 143.565 93.025 143.640 ;
        RECT 68.090 143.415 93.025 143.565 ;
        RECT 68.090 143.340 68.490 143.415 ;
        RECT 77.490 143.340 77.890 143.415 ;
        RECT 92.625 143.340 93.025 143.415 ;
        RECT 96.075 143.565 96.475 143.640 ;
        RECT 157.350 143.565 157.500 189.340 ;
        RECT 96.075 143.415 157.500 143.565 ;
        RECT 96.075 143.340 96.475 143.415 ;
        RECT 7.290 142.565 35.940 142.915 ;
        RECT 7.290 133.415 7.690 142.565 ;
        RECT 8.240 142.270 8.640 142.315 ;
        RECT 8.240 142.020 18.240 142.270 ;
        RECT 18.490 142.265 18.890 142.315 ;
        RECT 23.590 142.265 23.990 142.315 ;
        RECT 26.190 142.265 26.590 142.315 ;
        RECT 8.240 142.015 8.640 142.020 ;
        RECT 18.440 142.015 23.390 142.265 ;
        RECT 23.590 142.015 25.940 142.265 ;
        RECT 26.140 142.015 27.190 142.265 ;
        RECT 27.440 142.015 27.840 142.315 ;
        RECT 28.640 142.015 29.040 142.315 ;
        RECT 29.890 142.015 30.290 142.315 ;
        RECT 31.090 142.015 31.490 142.315 ;
        RECT 32.290 142.015 32.690 142.315 ;
        RECT 33.540 142.015 33.940 142.315 ;
        RECT 34.690 142.015 35.090 142.315 ;
        RECT 8.005 138.565 8.235 141.815 ;
        RECT 7.890 138.265 8.290 138.565 ;
        RECT 8.005 133.815 8.235 138.265 ;
        RECT 8.645 134.215 8.875 141.815 ;
        RECT 9.285 138.565 9.515 141.815 ;
        RECT 9.190 138.265 9.590 138.565 ;
        RECT 8.540 133.915 8.940 134.215 ;
        RECT 8.645 133.815 8.875 133.915 ;
        RECT 9.285 133.815 9.515 138.265 ;
        RECT 9.925 134.215 10.155 141.815 ;
        RECT 10.565 138.565 10.795 141.815 ;
        RECT 10.490 138.265 10.890 138.565 ;
        RECT 9.840 133.915 10.240 134.215 ;
        RECT 9.925 133.815 10.155 133.915 ;
        RECT 10.565 133.815 10.795 138.265 ;
        RECT 11.205 134.215 11.435 141.815 ;
        RECT 11.845 138.565 12.075 141.815 ;
        RECT 11.740 138.265 12.140 138.565 ;
        RECT 11.140 133.915 11.540 134.215 ;
        RECT 11.205 133.815 11.435 133.915 ;
        RECT 11.845 133.815 12.075 138.265 ;
        RECT 12.485 134.215 12.715 141.815 ;
        RECT 13.125 138.565 13.355 141.815 ;
        RECT 13.040 138.265 13.440 138.565 ;
        RECT 12.390 133.915 12.790 134.215 ;
        RECT 12.485 133.815 12.715 133.915 ;
        RECT 13.125 133.815 13.355 138.265 ;
        RECT 13.765 134.215 13.995 141.815 ;
        RECT 14.405 138.565 14.635 141.815 ;
        RECT 14.290 138.265 14.690 138.565 ;
        RECT 13.690 133.915 14.090 134.215 ;
        RECT 13.765 133.815 13.995 133.915 ;
        RECT 14.405 133.815 14.635 138.265 ;
        RECT 15.045 134.215 15.275 141.815 ;
        RECT 15.685 138.565 15.915 141.815 ;
        RECT 15.590 138.265 15.990 138.565 ;
        RECT 14.940 133.915 15.340 134.215 ;
        RECT 15.045 133.815 15.275 133.915 ;
        RECT 15.685 133.815 15.915 138.265 ;
        RECT 16.325 134.215 16.555 141.815 ;
        RECT 16.965 138.565 17.195 141.815 ;
        RECT 16.890 138.265 17.290 138.565 ;
        RECT 16.240 133.915 16.640 134.215 ;
        RECT 16.325 133.815 16.555 133.915 ;
        RECT 16.965 133.815 17.195 138.265 ;
        RECT 17.605 134.215 17.835 141.815 ;
        RECT 18.245 138.565 18.475 141.815 ;
        RECT 18.140 138.265 18.540 138.565 ;
        RECT 17.540 133.915 17.940 134.215 ;
        RECT 17.605 133.815 17.835 133.915 ;
        RECT 18.245 133.815 18.475 138.265 ;
        RECT 18.885 134.215 19.115 141.815 ;
        RECT 19.525 138.565 19.755 141.815 ;
        RECT 19.440 138.265 19.840 138.565 ;
        RECT 18.790 133.915 19.190 134.215 ;
        RECT 18.885 133.815 19.115 133.915 ;
        RECT 19.525 133.815 19.755 138.265 ;
        RECT 20.165 134.215 20.395 141.815 ;
        RECT 20.805 138.565 21.035 141.815 ;
        RECT 20.690 138.265 21.090 138.565 ;
        RECT 20.090 133.915 20.490 134.215 ;
        RECT 20.165 133.815 20.395 133.915 ;
        RECT 20.805 133.815 21.035 138.265 ;
        RECT 21.445 134.215 21.675 141.815 ;
        RECT 22.085 138.565 22.315 141.815 ;
        RECT 21.990 138.265 22.390 138.565 ;
        RECT 21.340 133.915 21.740 134.215 ;
        RECT 21.445 133.815 21.675 133.915 ;
        RECT 22.085 133.815 22.315 138.265 ;
        RECT 22.725 134.215 22.955 141.815 ;
        RECT 23.365 138.565 23.595 141.815 ;
        RECT 23.290 138.265 23.690 138.565 ;
        RECT 22.640 133.915 23.040 134.215 ;
        RECT 22.725 133.815 22.955 133.915 ;
        RECT 23.365 133.815 23.595 138.265 ;
        RECT 24.005 134.215 24.235 141.815 ;
        RECT 24.645 138.565 24.875 141.815 ;
        RECT 24.540 138.265 24.940 138.565 ;
        RECT 23.890 133.915 24.290 134.215 ;
        RECT 24.005 133.815 24.235 133.915 ;
        RECT 24.645 133.815 24.875 138.265 ;
        RECT 25.285 134.215 25.515 141.815 ;
        RECT 25.925 138.565 26.155 141.815 ;
        RECT 25.840 138.265 26.240 138.565 ;
        RECT 25.190 133.915 25.590 134.215 ;
        RECT 25.285 133.815 25.515 133.915 ;
        RECT 25.925 133.815 26.155 138.265 ;
        RECT 26.565 134.215 26.795 141.815 ;
        RECT 27.205 138.565 27.435 141.815 ;
        RECT 27.140 138.265 27.540 138.565 ;
        RECT 26.490 133.915 26.890 134.215 ;
        RECT 26.565 133.815 26.795 133.915 ;
        RECT 27.205 133.815 27.435 138.265 ;
        RECT 27.845 134.215 28.075 141.815 ;
        RECT 28.430 138.565 28.660 141.815 ;
        RECT 28.340 138.265 28.740 138.565 ;
        RECT 28.430 137.815 28.660 138.265 ;
        RECT 29.070 137.815 29.300 141.815 ;
        RECT 29.640 138.565 29.870 141.815 ;
        RECT 29.540 138.265 29.940 138.565 ;
        RECT 29.640 137.815 29.870 138.265 ;
        RECT 30.280 137.815 30.510 141.815 ;
        RECT 30.850 138.565 31.080 141.815 ;
        RECT 30.740 138.265 31.140 138.565 ;
        RECT 30.850 137.815 31.080 138.265 ;
        RECT 31.490 137.815 31.720 141.815 ;
        RECT 32.060 138.565 32.290 141.815 ;
        RECT 31.990 138.265 32.390 138.565 ;
        RECT 32.700 138.265 32.930 141.815 ;
        RECT 33.270 138.565 33.500 141.815 ;
        RECT 33.190 138.265 33.590 138.565 ;
        RECT 32.060 137.815 32.290 138.265 ;
        RECT 32.700 137.815 32.940 138.265 ;
        RECT 33.270 137.815 33.500 138.265 ;
        RECT 33.910 137.815 34.140 141.815 ;
        RECT 34.480 138.565 34.710 141.815 ;
        RECT 34.390 138.265 34.790 138.565 ;
        RECT 34.480 137.815 34.710 138.265 ;
        RECT 35.120 137.815 35.350 141.815 ;
        RECT 27.740 133.915 28.140 134.215 ;
        RECT 29.090 134.065 29.290 137.815 ;
        RECT 30.290 134.065 30.490 137.815 ;
        RECT 31.490 134.065 31.690 137.815 ;
        RECT 32.740 134.065 32.940 137.815 ;
        RECT 33.940 134.065 34.140 137.815 ;
        RECT 35.140 134.065 35.340 137.815 ;
        RECT 27.845 133.815 28.075 133.915 ;
        RECT 28.990 133.765 29.390 134.065 ;
        RECT 30.190 133.765 30.590 134.065 ;
        RECT 31.390 133.765 31.790 134.065 ;
        RECT 32.640 133.765 33.040 134.065 ;
        RECT 33.840 133.765 34.240 134.065 ;
        RECT 35.040 133.765 35.440 134.065 ;
        RECT 35.690 133.415 35.940 142.565 ;
        RECT 7.290 133.065 35.940 133.415 ;
        RECT 36.090 142.565 75.290 142.915 ;
        RECT 36.090 133.415 36.440 142.565 ;
        RECT 37.440 142.165 37.840 142.215 ;
        RECT 41.290 142.165 41.690 142.215 ;
        RECT 37.440 141.915 40.740 142.165 ;
        RECT 41.290 141.915 42.640 142.165 ;
        RECT 43.240 141.915 43.640 142.215 ;
        RECT 44.090 141.915 44.490 142.215 ;
        RECT 45.190 141.915 46.490 142.215 ;
        RECT 47.290 141.915 50.590 142.215 ;
        RECT 51.140 141.915 54.390 142.215 ;
        RECT 54.990 141.915 56.290 142.215 ;
        RECT 56.890 141.915 57.290 142.215 ;
        RECT 57.840 141.915 58.240 142.215 ;
        RECT 58.890 141.915 59.290 142.215 ;
        RECT 59.840 141.915 60.240 142.215 ;
        RECT 60.440 141.915 60.840 142.215 ;
        RECT 61.490 141.915 61.890 142.215 ;
        RECT 62.540 141.915 62.940 142.215 ;
        RECT 63.590 141.915 63.990 142.215 ;
        RECT 64.640 141.915 65.040 142.215 ;
        RECT 72.240 142.115 73.290 142.315 ;
        RECT 36.825 136.515 37.055 141.775 ;
        RECT 36.740 136.215 37.140 136.515 ;
        RECT 36.825 133.775 37.055 136.215 ;
        RECT 37.305 134.315 37.535 141.775 ;
        RECT 37.785 136.515 38.015 141.775 ;
        RECT 37.690 136.215 38.090 136.515 ;
        RECT 37.240 134.015 37.640 134.315 ;
        RECT 37.305 133.775 37.535 134.015 ;
        RECT 37.785 133.775 38.015 136.215 ;
        RECT 38.265 134.315 38.495 141.775 ;
        RECT 38.745 136.515 38.975 141.775 ;
        RECT 38.640 136.215 39.040 136.515 ;
        RECT 38.190 134.015 38.590 134.315 ;
        RECT 38.265 133.775 38.495 134.015 ;
        RECT 38.745 133.775 38.975 136.215 ;
        RECT 39.225 134.315 39.455 141.775 ;
        RECT 39.705 136.515 39.935 141.775 ;
        RECT 39.640 136.215 40.040 136.515 ;
        RECT 39.140 134.015 39.540 134.315 ;
        RECT 39.225 133.775 39.455 134.015 ;
        RECT 39.705 133.775 39.935 136.215 ;
        RECT 40.185 134.315 40.415 141.775 ;
        RECT 40.665 136.515 40.895 141.775 ;
        RECT 40.590 136.215 40.990 136.515 ;
        RECT 40.090 134.015 40.490 134.315 ;
        RECT 40.185 133.775 40.415 134.015 ;
        RECT 40.665 133.775 40.895 136.215 ;
        RECT 41.145 134.315 41.375 141.775 ;
        RECT 41.625 136.515 41.855 141.775 ;
        RECT 41.540 136.215 41.940 136.515 ;
        RECT 41.040 134.015 41.440 134.315 ;
        RECT 41.145 133.775 41.375 134.015 ;
        RECT 41.625 133.775 41.855 136.215 ;
        RECT 42.105 134.315 42.335 141.775 ;
        RECT 42.585 136.515 42.815 141.775 ;
        RECT 42.490 136.215 42.890 136.515 ;
        RECT 42.040 134.015 42.440 134.315 ;
        RECT 42.105 133.775 42.335 134.015 ;
        RECT 42.585 133.775 42.815 136.215 ;
        RECT 43.065 134.315 43.295 141.775 ;
        RECT 43.545 136.515 43.775 141.775 ;
        RECT 43.440 136.215 43.840 136.515 ;
        RECT 42.990 134.015 43.390 134.315 ;
        RECT 43.065 133.775 43.295 134.015 ;
        RECT 43.545 133.775 43.775 136.215 ;
        RECT 44.025 134.315 44.255 141.775 ;
        RECT 44.590 135.865 44.820 141.775 ;
        RECT 44.490 135.565 44.890 135.865 ;
        RECT 43.940 134.015 44.340 134.315 ;
        RECT 44.025 133.775 44.255 134.015 ;
        RECT 44.590 133.775 44.820 135.565 ;
        RECT 45.070 134.315 45.300 141.775 ;
        RECT 45.550 135.865 45.780 141.775 ;
        RECT 45.440 135.565 45.840 135.865 ;
        RECT 44.990 134.015 45.390 134.315 ;
        RECT 45.070 133.775 45.300 134.015 ;
        RECT 45.550 133.775 45.780 135.565 ;
        RECT 46.030 134.315 46.260 141.775 ;
        RECT 46.670 141.615 46.900 141.775 ;
        RECT 46.590 141.315 46.990 141.615 ;
        RECT 45.940 134.015 46.340 134.315 ;
        RECT 46.030 133.775 46.260 134.015 ;
        RECT 46.670 133.775 46.900 141.315 ;
        RECT 47.150 140.615 47.380 141.775 ;
        RECT 47.630 141.615 47.860 141.775 ;
        RECT 47.540 141.315 47.940 141.615 ;
        RECT 47.090 140.315 47.490 140.615 ;
        RECT 47.150 133.775 47.380 140.315 ;
        RECT 47.630 133.775 47.860 141.315 ;
        RECT 48.110 140.615 48.340 141.775 ;
        RECT 48.590 141.615 48.820 141.775 ;
        RECT 48.490 141.315 48.890 141.615 ;
        RECT 48.040 140.315 48.440 140.615 ;
        RECT 48.110 133.775 48.340 140.315 ;
        RECT 48.590 133.775 48.820 141.315 ;
        RECT 49.070 140.615 49.300 141.775 ;
        RECT 49.550 141.615 49.780 141.775 ;
        RECT 49.440 141.315 49.840 141.615 ;
        RECT 48.990 140.315 49.390 140.615 ;
        RECT 49.070 133.775 49.300 140.315 ;
        RECT 49.550 133.775 49.780 141.315 ;
        RECT 50.030 140.615 50.260 141.775 ;
        RECT 50.510 141.615 50.740 141.775 ;
        RECT 50.440 141.315 50.840 141.615 ;
        RECT 49.940 140.315 50.340 140.615 ;
        RECT 50.030 133.775 50.260 140.315 ;
        RECT 50.510 133.775 50.740 141.315 ;
        RECT 50.990 134.165 51.220 141.775 ;
        RECT 51.470 141.615 51.700 141.775 ;
        RECT 51.390 141.315 51.790 141.615 ;
        RECT 50.890 133.865 51.290 134.165 ;
        RECT 50.990 133.775 51.220 133.865 ;
        RECT 51.470 133.775 51.700 141.315 ;
        RECT 51.950 134.165 52.180 141.775 ;
        RECT 52.430 141.615 52.660 141.775 ;
        RECT 52.340 141.315 52.740 141.615 ;
        RECT 51.890 133.865 52.290 134.165 ;
        RECT 51.950 133.775 52.180 133.865 ;
        RECT 52.430 133.775 52.660 141.315 ;
        RECT 52.910 134.165 53.140 141.775 ;
        RECT 53.390 141.615 53.620 141.775 ;
        RECT 53.290 141.315 53.690 141.615 ;
        RECT 52.840 133.865 53.240 134.165 ;
        RECT 52.910 133.775 53.140 133.865 ;
        RECT 53.390 133.775 53.620 141.315 ;
        RECT 53.870 134.165 54.100 141.775 ;
        RECT 54.350 141.615 54.580 141.775 ;
        RECT 54.290 141.315 54.690 141.615 ;
        RECT 53.790 133.865 54.190 134.165 ;
        RECT 53.870 133.775 54.100 133.865 ;
        RECT 54.350 133.775 54.580 141.315 ;
        RECT 54.830 134.165 55.060 141.775 ;
        RECT 55.310 141.615 55.540 141.775 ;
        RECT 55.240 141.315 55.640 141.615 ;
        RECT 54.740 133.865 55.140 134.165 ;
        RECT 54.830 133.775 55.060 133.865 ;
        RECT 55.310 133.775 55.540 141.315 ;
        RECT 55.790 134.165 56.020 141.775 ;
        RECT 56.270 141.615 56.500 141.775 ;
        RECT 56.190 141.315 56.590 141.615 ;
        RECT 55.690 133.865 56.090 134.165 ;
        RECT 55.790 133.775 56.020 133.865 ;
        RECT 56.270 133.775 56.500 141.315 ;
        RECT 56.750 134.165 56.980 141.775 ;
        RECT 57.230 141.615 57.460 141.775 ;
        RECT 57.140 141.315 57.540 141.615 ;
        RECT 56.690 133.865 57.090 134.165 ;
        RECT 56.750 133.775 56.980 133.865 ;
        RECT 57.230 133.775 57.460 141.315 ;
        RECT 57.710 134.165 57.940 141.775 ;
        RECT 58.270 141.115 58.500 141.775 ;
        RECT 58.190 140.815 58.590 141.115 ;
        RECT 58.270 139.775 58.500 140.815 ;
        RECT 58.750 140.265 58.980 141.775 ;
        RECT 59.230 141.115 59.460 141.775 ;
        RECT 59.140 140.815 59.540 141.115 ;
        RECT 58.690 139.965 59.090 140.265 ;
        RECT 58.750 139.775 58.980 139.965 ;
        RECT 59.230 139.775 59.460 140.815 ;
        RECT 59.710 140.265 59.940 141.775 ;
        RECT 60.270 141.115 60.500 141.775 ;
        RECT 60.190 140.815 60.590 141.115 ;
        RECT 59.640 139.965 60.040 140.265 ;
        RECT 59.710 139.775 59.940 139.965 ;
        RECT 60.270 139.775 60.500 140.815 ;
        RECT 60.750 140.265 60.980 141.775 ;
        RECT 61.320 141.115 61.550 141.775 ;
        RECT 61.240 140.815 61.640 141.115 ;
        RECT 60.690 139.965 61.090 140.265 ;
        RECT 60.750 139.775 60.980 139.965 ;
        RECT 61.320 139.775 61.550 140.815 ;
        RECT 61.800 140.265 62.030 141.775 ;
        RECT 62.370 141.115 62.600 141.775 ;
        RECT 62.290 140.815 62.690 141.115 ;
        RECT 61.740 139.965 62.140 140.265 ;
        RECT 61.800 139.775 62.030 139.965 ;
        RECT 62.370 139.775 62.600 140.815 ;
        RECT 62.850 140.265 63.080 141.775 ;
        RECT 63.420 141.115 63.650 141.775 ;
        RECT 63.340 140.815 63.740 141.115 ;
        RECT 62.790 139.965 63.190 140.265 ;
        RECT 62.850 139.775 63.080 139.965 ;
        RECT 63.420 139.775 63.650 140.815 ;
        RECT 63.900 140.315 64.130 141.775 ;
        RECT 64.470 141.115 64.700 141.775 ;
        RECT 64.390 140.815 64.790 141.115 ;
        RECT 63.840 140.015 64.240 140.315 ;
        RECT 63.900 139.775 64.130 140.015 ;
        RECT 64.470 139.775 64.700 140.815 ;
        RECT 64.950 140.315 65.180 141.775 ;
        RECT 64.890 140.015 65.290 140.315 ;
        RECT 72.240 140.265 72.490 142.115 ;
        RECT 72.970 142.070 73.260 142.115 ;
        RECT 72.760 141.565 72.990 141.910 ;
        RECT 72.640 141.265 73.040 141.565 ;
        RECT 73.240 141.265 73.470 141.910 ;
        RECT 74.440 141.265 74.840 141.365 ;
        RECT 72.760 140.910 72.990 141.265 ;
        RECT 73.240 141.115 74.840 141.265 ;
        RECT 73.240 140.910 73.470 141.115 ;
        RECT 74.440 141.065 74.840 141.115 ;
        RECT 72.970 140.265 73.260 140.285 ;
        RECT 72.240 140.065 73.290 140.265 ;
        RECT 64.950 139.775 65.180 140.015 ;
        RECT 64.140 139.515 64.540 139.565 ;
        RECT 72.240 139.515 72.490 140.065 ;
        RECT 72.970 140.055 73.260 140.065 ;
        RECT 72.760 139.515 72.990 139.895 ;
        RECT 64.140 139.315 72.490 139.515 ;
        RECT 64.140 139.265 64.540 139.315 ;
        RECT 68.090 139.115 68.490 139.165 ;
        RECT 58.940 138.915 68.490 139.115 ;
        RECT 58.940 138.815 59.340 138.915 ;
        RECT 68.090 138.865 68.490 138.915 ;
        RECT 59.890 138.715 60.290 138.765 ;
        RECT 67.290 138.715 67.690 138.765 ;
        RECT 59.890 138.515 67.690 138.715 ;
        RECT 59.890 138.465 60.290 138.515 ;
        RECT 67.290 138.465 67.690 138.515 ;
        RECT 60.440 138.315 60.840 138.365 ;
        RECT 66.490 138.315 66.890 138.365 ;
        RECT 60.440 138.115 66.890 138.315 ;
        RECT 60.440 138.065 60.840 138.115 ;
        RECT 66.490 138.065 66.890 138.115 ;
        RECT 72.240 138.115 72.490 139.315 ;
        RECT 72.640 139.215 73.040 139.515 ;
        RECT 73.240 139.265 73.470 139.895 ;
        RECT 74.040 139.265 74.440 139.365 ;
        RECT 72.760 138.895 72.990 139.215 ;
        RECT 73.240 139.115 74.440 139.265 ;
        RECT 73.240 138.895 73.470 139.115 ;
        RECT 74.040 139.065 74.440 139.115 ;
        RECT 72.980 138.115 73.270 138.120 ;
        RECT 61.490 137.915 61.890 137.965 ;
        RECT 67.690 137.915 68.090 137.965 ;
        RECT 61.490 137.715 68.090 137.915 ;
        RECT 61.490 137.665 61.890 137.715 ;
        RECT 67.690 137.665 68.090 137.715 ;
        RECT 72.240 137.915 73.290 138.115 ;
        RECT 62.540 137.515 62.940 137.565 ;
        RECT 66.890 137.515 67.290 137.565 ;
        RECT 62.540 137.315 67.290 137.515 ;
        RECT 62.540 137.265 62.940 137.315 ;
        RECT 66.890 137.265 67.290 137.315 ;
        RECT 63.590 137.115 63.990 137.165 ;
        RECT 66.090 137.115 66.490 137.165 ;
        RECT 63.590 136.915 66.490 137.115 ;
        RECT 63.590 136.865 63.990 136.915 ;
        RECT 66.090 136.865 66.490 136.915 ;
        RECT 64.640 136.715 65.040 136.765 ;
        RECT 65.290 136.715 65.690 136.765 ;
        RECT 64.640 136.515 65.690 136.715 ;
        RECT 64.640 136.465 65.040 136.515 ;
        RECT 65.290 136.465 65.690 136.515 ;
        RECT 72.240 136.215 72.490 137.915 ;
        RECT 72.980 137.890 73.270 137.915 ;
        RECT 72.770 137.365 73.000 137.730 ;
        RECT 72.640 137.065 73.040 137.365 ;
        RECT 72.770 136.730 73.000 137.065 ;
        RECT 73.250 137.015 73.480 137.730 ;
        RECT 73.640 137.015 74.040 137.115 ;
        RECT 73.250 136.865 74.040 137.015 ;
        RECT 73.250 136.730 73.480 136.865 ;
        RECT 73.640 136.815 74.040 136.865 ;
        RECT 58.940 135.915 59.340 136.215 ;
        RECT 59.890 135.915 60.290 136.215 ;
        RECT 60.440 135.915 60.840 136.215 ;
        RECT 61.490 135.915 61.890 136.215 ;
        RECT 62.540 135.915 62.940 136.215 ;
        RECT 63.590 135.915 63.990 136.215 ;
        RECT 64.640 135.915 65.040 136.215 ;
        RECT 65.690 135.915 66.090 136.215 ;
        RECT 67.240 135.965 73.290 136.215 ;
        RECT 67.260 135.940 67.550 135.965 ;
        RECT 68.220 135.940 68.510 135.965 ;
        RECT 68.780 135.940 69.070 135.965 ;
        RECT 69.830 135.940 70.120 135.965 ;
        RECT 70.880 135.940 71.170 135.965 ;
        RECT 71.930 135.940 72.220 135.965 ;
        RECT 72.980 135.940 73.270 135.965 ;
        RECT 58.270 135.665 58.500 135.775 ;
        RECT 58.190 135.365 58.590 135.665 ;
        RECT 57.640 133.865 58.040 134.165 ;
        RECT 57.710 133.775 57.940 133.865 ;
        RECT 58.270 133.775 58.500 135.365 ;
        RECT 58.750 134.365 58.980 135.775 ;
        RECT 59.230 135.665 59.460 135.775 ;
        RECT 59.140 135.365 59.540 135.665 ;
        RECT 58.690 134.065 59.090 134.365 ;
        RECT 58.750 133.775 58.980 134.065 ;
        RECT 59.230 133.775 59.460 135.365 ;
        RECT 59.710 134.365 59.940 135.775 ;
        RECT 60.270 135.665 60.500 135.775 ;
        RECT 60.190 135.365 60.590 135.665 ;
        RECT 59.640 134.065 60.040 134.365 ;
        RECT 59.710 133.775 59.940 134.065 ;
        RECT 60.270 133.775 60.500 135.365 ;
        RECT 60.750 134.365 60.980 135.775 ;
        RECT 61.320 135.665 61.550 135.775 ;
        RECT 61.240 135.365 61.640 135.665 ;
        RECT 60.690 134.065 61.090 134.365 ;
        RECT 60.750 133.775 60.980 134.065 ;
        RECT 61.320 133.775 61.550 135.365 ;
        RECT 61.800 134.365 62.030 135.775 ;
        RECT 62.370 135.665 62.600 135.775 ;
        RECT 62.290 135.365 62.690 135.665 ;
        RECT 61.740 134.065 62.140 134.365 ;
        RECT 61.800 133.775 62.030 134.065 ;
        RECT 62.370 133.775 62.600 135.365 ;
        RECT 62.850 134.365 63.080 135.775 ;
        RECT 63.420 135.665 63.650 135.775 ;
        RECT 63.340 135.365 63.740 135.665 ;
        RECT 62.790 134.065 63.190 134.365 ;
        RECT 62.850 133.775 63.080 134.065 ;
        RECT 63.420 133.775 63.650 135.365 ;
        RECT 63.900 134.365 64.130 135.775 ;
        RECT 64.470 135.665 64.700 135.775 ;
        RECT 64.390 135.365 64.790 135.665 ;
        RECT 63.840 134.065 64.240 134.365 ;
        RECT 63.900 133.775 64.130 134.065 ;
        RECT 64.470 133.775 64.700 135.365 ;
        RECT 64.950 134.365 65.180 135.775 ;
        RECT 65.520 135.665 65.750 135.775 ;
        RECT 65.440 135.365 65.840 135.665 ;
        RECT 64.890 134.065 65.290 134.365 ;
        RECT 64.950 133.775 65.180 134.065 ;
        RECT 65.520 133.775 65.750 135.365 ;
        RECT 66.000 134.365 66.230 135.775 ;
        RECT 66.570 135.665 66.800 135.780 ;
        RECT 66.490 135.365 66.890 135.665 ;
        RECT 65.940 134.065 66.340 134.365 ;
        RECT 66.000 133.775 66.230 134.065 ;
        RECT 66.570 133.780 66.800 135.365 ;
        RECT 67.050 134.215 67.280 135.780 ;
        RECT 67.530 135.665 67.760 135.780 ;
        RECT 67.440 135.365 67.840 135.665 ;
        RECT 66.990 133.915 67.390 134.215 ;
        RECT 67.050 133.780 67.280 133.915 ;
        RECT 67.530 133.780 67.760 135.365 ;
        RECT 68.010 134.215 68.240 135.780 ;
        RECT 68.570 135.115 68.800 135.780 ;
        RECT 69.050 135.665 69.280 135.780 ;
        RECT 68.990 135.365 69.390 135.665 ;
        RECT 68.490 134.815 68.890 135.115 ;
        RECT 68.570 134.780 68.800 134.815 ;
        RECT 69.050 134.780 69.280 135.365 ;
        RECT 69.620 135.115 69.850 135.780 ;
        RECT 70.100 135.665 70.330 135.780 ;
        RECT 70.040 135.365 70.440 135.665 ;
        RECT 69.540 134.815 69.940 135.115 ;
        RECT 69.620 134.780 69.850 134.815 ;
        RECT 70.100 134.780 70.330 135.365 ;
        RECT 70.670 135.115 70.900 135.780 ;
        RECT 71.150 135.665 71.380 135.780 ;
        RECT 71.090 135.365 71.490 135.665 ;
        RECT 70.590 134.815 70.990 135.115 ;
        RECT 70.670 134.780 70.900 134.815 ;
        RECT 71.150 134.780 71.380 135.365 ;
        RECT 71.720 135.115 71.950 135.780 ;
        RECT 72.200 135.665 72.430 135.780 ;
        RECT 72.140 135.365 72.540 135.665 ;
        RECT 71.640 134.815 72.040 135.115 ;
        RECT 71.720 134.780 71.950 134.815 ;
        RECT 72.200 134.780 72.430 135.365 ;
        RECT 72.770 135.115 73.000 135.780 ;
        RECT 73.250 135.665 73.480 135.780 ;
        RECT 73.190 135.365 73.590 135.665 ;
        RECT 72.690 134.815 73.090 135.115 ;
        RECT 72.770 134.780 73.000 134.815 ;
        RECT 73.250 134.780 73.480 135.365 ;
        RECT 67.940 133.915 68.340 134.215 ;
        RECT 68.010 133.780 68.240 133.915 ;
        RECT 74.990 133.415 75.290 142.565 ;
        RECT 36.090 133.065 75.290 133.415 ;
        RECT 85.825 142.565 125.025 142.915 ;
        RECT 85.825 133.415 86.125 142.565 ;
        RECT 87.825 142.115 88.875 142.315 ;
        RECT 87.855 142.070 88.145 142.115 ;
        RECT 86.275 141.265 86.675 141.365 ;
        RECT 87.645 141.265 87.875 141.910 ;
        RECT 88.125 141.565 88.355 141.910 ;
        RECT 88.075 141.265 88.475 141.565 ;
        RECT 86.275 141.115 87.875 141.265 ;
        RECT 86.275 141.065 86.675 141.115 ;
        RECT 87.645 140.910 87.875 141.115 ;
        RECT 88.125 140.910 88.355 141.265 ;
        RECT 87.855 140.265 88.145 140.285 ;
        RECT 88.625 140.265 88.875 142.115 ;
        RECT 96.075 141.915 96.475 142.215 ;
        RECT 97.125 141.915 97.525 142.215 ;
        RECT 98.175 141.915 98.575 142.215 ;
        RECT 99.225 141.915 99.625 142.215 ;
        RECT 100.275 141.915 100.675 142.215 ;
        RECT 100.875 141.915 101.275 142.215 ;
        RECT 101.825 141.915 102.225 142.215 ;
        RECT 102.875 141.915 103.275 142.215 ;
        RECT 103.825 141.915 104.225 142.215 ;
        RECT 104.825 141.915 106.125 142.215 ;
        RECT 106.725 141.915 109.975 142.215 ;
        RECT 110.525 141.915 113.825 142.215 ;
        RECT 114.625 141.915 115.925 142.215 ;
        RECT 116.625 141.915 117.025 142.215 ;
        RECT 117.475 141.915 117.875 142.215 ;
        RECT 119.425 142.165 119.825 142.215 ;
        RECT 123.275 142.165 123.675 142.215 ;
        RECT 118.475 141.915 119.825 142.165 ;
        RECT 120.375 141.915 123.675 142.165 ;
        RECT 95.935 140.315 96.165 141.775 ;
        RECT 96.415 141.115 96.645 141.775 ;
        RECT 96.325 140.815 96.725 141.115 ;
        RECT 87.825 140.065 88.875 140.265 ;
        RECT 87.855 140.055 88.145 140.065 ;
        RECT 86.675 139.265 87.075 139.365 ;
        RECT 87.645 139.265 87.875 139.895 ;
        RECT 88.125 139.515 88.355 139.895 ;
        RECT 88.625 139.515 88.875 140.065 ;
        RECT 95.825 140.015 96.225 140.315 ;
        RECT 95.935 139.775 96.165 140.015 ;
        RECT 96.415 139.775 96.645 140.815 ;
        RECT 96.985 140.315 97.215 141.775 ;
        RECT 97.465 141.115 97.695 141.775 ;
        RECT 97.375 140.815 97.775 141.115 ;
        RECT 96.875 140.015 97.275 140.315 ;
        RECT 96.985 139.775 97.215 140.015 ;
        RECT 97.465 139.775 97.695 140.815 ;
        RECT 98.035 140.265 98.265 141.775 ;
        RECT 98.515 141.115 98.745 141.775 ;
        RECT 98.425 140.815 98.825 141.115 ;
        RECT 97.925 139.965 98.325 140.265 ;
        RECT 98.035 139.775 98.265 139.965 ;
        RECT 98.515 139.775 98.745 140.815 ;
        RECT 99.085 140.265 99.315 141.775 ;
        RECT 99.565 141.115 99.795 141.775 ;
        RECT 99.475 140.815 99.875 141.115 ;
        RECT 98.975 139.965 99.375 140.265 ;
        RECT 99.085 139.775 99.315 139.965 ;
        RECT 99.565 139.775 99.795 140.815 ;
        RECT 100.135 140.265 100.365 141.775 ;
        RECT 100.615 141.115 100.845 141.775 ;
        RECT 100.525 140.815 100.925 141.115 ;
        RECT 100.025 139.965 100.425 140.265 ;
        RECT 100.135 139.775 100.365 139.965 ;
        RECT 100.615 139.775 100.845 140.815 ;
        RECT 101.175 140.265 101.405 141.775 ;
        RECT 101.655 141.115 101.885 141.775 ;
        RECT 101.575 140.815 101.975 141.115 ;
        RECT 101.075 139.965 101.475 140.265 ;
        RECT 101.175 139.775 101.405 139.965 ;
        RECT 101.655 139.775 101.885 140.815 ;
        RECT 102.135 140.265 102.365 141.775 ;
        RECT 102.615 141.115 102.845 141.775 ;
        RECT 102.525 140.815 102.925 141.115 ;
        RECT 102.025 139.965 102.425 140.265 ;
        RECT 102.135 139.775 102.365 139.965 ;
        RECT 102.615 139.775 102.845 140.815 ;
        RECT 96.575 139.515 96.975 139.565 ;
        RECT 86.675 139.115 87.875 139.265 ;
        RECT 88.075 139.215 88.475 139.515 ;
        RECT 88.625 139.315 96.975 139.515 ;
        RECT 86.675 139.065 87.075 139.115 ;
        RECT 87.645 138.895 87.875 139.115 ;
        RECT 88.125 138.895 88.355 139.215 ;
        RECT 87.845 138.115 88.135 138.120 ;
        RECT 88.625 138.115 88.875 139.315 ;
        RECT 96.575 139.265 96.975 139.315 ;
        RECT 92.625 139.115 93.025 139.165 ;
        RECT 92.625 138.915 102.175 139.115 ;
        RECT 92.625 138.865 93.025 138.915 ;
        RECT 101.775 138.815 102.175 138.915 ;
        RECT 93.425 138.715 93.825 138.765 ;
        RECT 100.825 138.715 101.225 138.765 ;
        RECT 93.425 138.515 101.225 138.715 ;
        RECT 93.425 138.465 93.825 138.515 ;
        RECT 100.825 138.465 101.225 138.515 ;
        RECT 87.825 137.915 88.875 138.115 ;
        RECT 94.225 138.315 94.625 138.365 ;
        RECT 100.275 138.315 100.675 138.365 ;
        RECT 94.225 138.115 100.675 138.315 ;
        RECT 94.225 138.065 94.625 138.115 ;
        RECT 100.275 138.065 100.675 138.115 ;
        RECT 87.845 137.890 88.135 137.915 ;
        RECT 87.075 137.015 87.475 137.115 ;
        RECT 87.635 137.015 87.865 137.730 ;
        RECT 88.115 137.365 88.345 137.730 ;
        RECT 88.075 137.065 88.475 137.365 ;
        RECT 87.075 136.865 87.865 137.015 ;
        RECT 87.075 136.815 87.475 136.865 ;
        RECT 87.635 136.730 87.865 136.865 ;
        RECT 88.115 136.730 88.345 137.065 ;
        RECT 88.625 136.215 88.875 137.915 ;
        RECT 93.025 137.915 93.425 137.965 ;
        RECT 99.225 137.915 99.625 137.965 ;
        RECT 93.025 137.715 99.625 137.915 ;
        RECT 93.025 137.665 93.425 137.715 ;
        RECT 99.225 137.665 99.625 137.715 ;
        RECT 93.825 137.515 94.225 137.565 ;
        RECT 98.175 137.515 98.575 137.565 ;
        RECT 93.825 137.315 98.575 137.515 ;
        RECT 93.825 137.265 94.225 137.315 ;
        RECT 98.175 137.265 98.575 137.315 ;
        RECT 94.625 137.115 95.025 137.165 ;
        RECT 97.125 137.115 97.525 137.165 ;
        RECT 94.625 136.915 97.525 137.115 ;
        RECT 94.625 136.865 95.025 136.915 ;
        RECT 97.125 136.865 97.525 136.915 ;
        RECT 95.425 136.715 95.825 136.765 ;
        RECT 96.075 136.715 96.475 136.765 ;
        RECT 95.425 136.515 96.475 136.715 ;
        RECT 95.425 136.465 95.825 136.515 ;
        RECT 96.075 136.465 96.475 136.515 ;
        RECT 87.825 135.965 93.875 136.215 ;
        RECT 87.845 135.940 88.135 135.965 ;
        RECT 88.895 135.940 89.185 135.965 ;
        RECT 89.945 135.940 90.235 135.965 ;
        RECT 90.995 135.940 91.285 135.965 ;
        RECT 92.045 135.940 92.335 135.965 ;
        RECT 92.605 135.940 92.895 135.965 ;
        RECT 93.565 135.940 93.855 135.965 ;
        RECT 95.025 135.915 95.425 136.215 ;
        RECT 96.075 135.915 96.475 136.215 ;
        RECT 97.125 135.915 97.525 136.215 ;
        RECT 98.175 135.915 98.575 136.215 ;
        RECT 99.225 135.915 99.625 136.215 ;
        RECT 100.275 135.915 100.675 136.215 ;
        RECT 100.825 135.915 101.225 136.215 ;
        RECT 101.775 135.915 102.175 136.215 ;
        RECT 87.635 135.665 87.865 135.780 ;
        RECT 87.525 135.365 87.925 135.665 ;
        RECT 87.635 134.780 87.865 135.365 ;
        RECT 88.115 135.115 88.345 135.780 ;
        RECT 88.685 135.665 88.915 135.780 ;
        RECT 88.575 135.365 88.975 135.665 ;
        RECT 88.025 134.815 88.425 135.115 ;
        RECT 88.115 134.780 88.345 134.815 ;
        RECT 88.685 134.780 88.915 135.365 ;
        RECT 89.165 135.115 89.395 135.780 ;
        RECT 89.735 135.665 89.965 135.780 ;
        RECT 89.625 135.365 90.025 135.665 ;
        RECT 89.075 134.815 89.475 135.115 ;
        RECT 89.165 134.780 89.395 134.815 ;
        RECT 89.735 134.780 89.965 135.365 ;
        RECT 90.215 135.115 90.445 135.780 ;
        RECT 90.785 135.665 91.015 135.780 ;
        RECT 90.675 135.365 91.075 135.665 ;
        RECT 90.125 134.815 90.525 135.115 ;
        RECT 90.215 134.780 90.445 134.815 ;
        RECT 90.785 134.780 91.015 135.365 ;
        RECT 91.265 135.115 91.495 135.780 ;
        RECT 91.835 135.665 92.065 135.780 ;
        RECT 91.725 135.365 92.125 135.665 ;
        RECT 91.175 134.815 91.575 135.115 ;
        RECT 91.265 134.780 91.495 134.815 ;
        RECT 91.835 134.780 92.065 135.365 ;
        RECT 92.315 135.115 92.545 135.780 ;
        RECT 92.225 134.815 92.625 135.115 ;
        RECT 92.315 134.780 92.545 134.815 ;
        RECT 92.875 134.215 93.105 135.780 ;
        RECT 93.355 135.665 93.585 135.780 ;
        RECT 93.275 135.365 93.675 135.665 ;
        RECT 92.775 133.915 93.175 134.215 ;
        RECT 92.875 133.780 93.105 133.915 ;
        RECT 93.355 133.780 93.585 135.365 ;
        RECT 93.835 134.215 94.065 135.780 ;
        RECT 94.315 135.665 94.545 135.780 ;
        RECT 94.225 135.365 94.625 135.665 ;
        RECT 93.725 133.915 94.125 134.215 ;
        RECT 93.835 133.780 94.065 133.915 ;
        RECT 94.315 133.780 94.545 135.365 ;
        RECT 94.885 134.365 95.115 135.775 ;
        RECT 95.365 135.665 95.595 135.775 ;
        RECT 95.275 135.365 95.675 135.665 ;
        RECT 94.775 134.065 95.175 134.365 ;
        RECT 94.885 133.775 95.115 134.065 ;
        RECT 95.365 133.775 95.595 135.365 ;
        RECT 95.935 134.365 96.165 135.775 ;
        RECT 96.415 135.665 96.645 135.775 ;
        RECT 96.325 135.365 96.725 135.665 ;
        RECT 95.825 134.065 96.225 134.365 ;
        RECT 95.935 133.775 96.165 134.065 ;
        RECT 96.415 133.775 96.645 135.365 ;
        RECT 96.985 134.365 97.215 135.775 ;
        RECT 97.465 135.665 97.695 135.775 ;
        RECT 97.375 135.365 97.775 135.665 ;
        RECT 96.875 134.065 97.275 134.365 ;
        RECT 96.985 133.775 97.215 134.065 ;
        RECT 97.465 133.775 97.695 135.365 ;
        RECT 98.035 134.365 98.265 135.775 ;
        RECT 98.515 135.665 98.745 135.775 ;
        RECT 98.425 135.365 98.825 135.665 ;
        RECT 97.925 134.065 98.325 134.365 ;
        RECT 98.035 133.775 98.265 134.065 ;
        RECT 98.515 133.775 98.745 135.365 ;
        RECT 99.085 134.365 99.315 135.775 ;
        RECT 99.565 135.665 99.795 135.775 ;
        RECT 99.475 135.365 99.875 135.665 ;
        RECT 98.975 134.065 99.375 134.365 ;
        RECT 99.085 133.775 99.315 134.065 ;
        RECT 99.565 133.775 99.795 135.365 ;
        RECT 100.135 134.365 100.365 135.775 ;
        RECT 100.615 135.665 100.845 135.775 ;
        RECT 100.525 135.365 100.925 135.665 ;
        RECT 100.025 134.065 100.425 134.365 ;
        RECT 100.135 133.775 100.365 134.065 ;
        RECT 100.615 133.775 100.845 135.365 ;
        RECT 101.175 134.365 101.405 135.775 ;
        RECT 101.655 135.665 101.885 135.775 ;
        RECT 101.575 135.365 101.975 135.665 ;
        RECT 101.075 134.065 101.475 134.365 ;
        RECT 101.175 133.775 101.405 134.065 ;
        RECT 101.655 133.775 101.885 135.365 ;
        RECT 102.135 134.365 102.365 135.775 ;
        RECT 102.615 135.665 102.845 135.775 ;
        RECT 102.525 135.365 102.925 135.665 ;
        RECT 102.025 134.065 102.425 134.365 ;
        RECT 102.135 133.775 102.365 134.065 ;
        RECT 102.615 133.775 102.845 135.365 ;
        RECT 103.175 134.165 103.405 141.775 ;
        RECT 103.655 141.615 103.885 141.775 ;
        RECT 103.575 141.315 103.975 141.615 ;
        RECT 103.075 133.865 103.475 134.165 ;
        RECT 103.175 133.775 103.405 133.865 ;
        RECT 103.655 133.775 103.885 141.315 ;
        RECT 104.135 134.165 104.365 141.775 ;
        RECT 104.615 141.615 104.845 141.775 ;
        RECT 104.525 141.315 104.925 141.615 ;
        RECT 104.025 133.865 104.425 134.165 ;
        RECT 104.135 133.775 104.365 133.865 ;
        RECT 104.615 133.775 104.845 141.315 ;
        RECT 105.095 134.165 105.325 141.775 ;
        RECT 105.575 141.615 105.805 141.775 ;
        RECT 105.475 141.315 105.875 141.615 ;
        RECT 105.025 133.865 105.425 134.165 ;
        RECT 105.095 133.775 105.325 133.865 ;
        RECT 105.575 133.775 105.805 141.315 ;
        RECT 106.055 134.165 106.285 141.775 ;
        RECT 106.535 141.615 106.765 141.775 ;
        RECT 106.425 141.315 106.825 141.615 ;
        RECT 105.975 133.865 106.375 134.165 ;
        RECT 106.055 133.775 106.285 133.865 ;
        RECT 106.535 133.775 106.765 141.315 ;
        RECT 107.015 134.165 107.245 141.775 ;
        RECT 107.495 141.615 107.725 141.775 ;
        RECT 107.425 141.315 107.825 141.615 ;
        RECT 106.925 133.865 107.325 134.165 ;
        RECT 107.015 133.775 107.245 133.865 ;
        RECT 107.495 133.775 107.725 141.315 ;
        RECT 107.975 134.165 108.205 141.775 ;
        RECT 108.455 141.615 108.685 141.775 ;
        RECT 108.375 141.315 108.775 141.615 ;
        RECT 107.875 133.865 108.275 134.165 ;
        RECT 107.975 133.775 108.205 133.865 ;
        RECT 108.455 133.775 108.685 141.315 ;
        RECT 108.935 134.165 109.165 141.775 ;
        RECT 109.415 141.615 109.645 141.775 ;
        RECT 109.325 141.315 109.725 141.615 ;
        RECT 108.825 133.865 109.225 134.165 ;
        RECT 108.935 133.775 109.165 133.865 ;
        RECT 109.415 133.775 109.645 141.315 ;
        RECT 109.895 134.165 110.125 141.775 ;
        RECT 110.375 141.615 110.605 141.775 ;
        RECT 110.275 141.315 110.675 141.615 ;
        RECT 109.825 133.865 110.225 134.165 ;
        RECT 109.895 133.775 110.125 133.865 ;
        RECT 110.375 133.775 110.605 141.315 ;
        RECT 110.855 140.615 111.085 141.775 ;
        RECT 111.335 141.615 111.565 141.775 ;
        RECT 111.275 141.315 111.675 141.615 ;
        RECT 110.775 140.315 111.175 140.615 ;
        RECT 110.855 133.775 111.085 140.315 ;
        RECT 111.335 133.775 111.565 141.315 ;
        RECT 111.815 140.615 112.045 141.775 ;
        RECT 112.295 141.615 112.525 141.775 ;
        RECT 112.225 141.315 112.625 141.615 ;
        RECT 111.725 140.315 112.125 140.615 ;
        RECT 111.815 133.775 112.045 140.315 ;
        RECT 112.295 133.775 112.525 141.315 ;
        RECT 112.775 140.615 113.005 141.775 ;
        RECT 113.255 141.615 113.485 141.775 ;
        RECT 113.175 141.315 113.575 141.615 ;
        RECT 112.675 140.315 113.075 140.615 ;
        RECT 112.775 133.775 113.005 140.315 ;
        RECT 113.255 133.775 113.485 141.315 ;
        RECT 113.735 140.615 113.965 141.775 ;
        RECT 114.215 141.615 114.445 141.775 ;
        RECT 114.125 141.315 114.525 141.615 ;
        RECT 113.625 140.315 114.025 140.615 ;
        RECT 113.735 133.775 113.965 140.315 ;
        RECT 114.215 133.775 114.445 141.315 ;
        RECT 114.855 134.315 115.085 141.775 ;
        RECT 115.335 135.865 115.565 141.775 ;
        RECT 115.275 135.565 115.675 135.865 ;
        RECT 114.775 134.015 115.175 134.315 ;
        RECT 114.855 133.775 115.085 134.015 ;
        RECT 115.335 133.775 115.565 135.565 ;
        RECT 115.815 134.315 116.045 141.775 ;
        RECT 116.295 135.865 116.525 141.775 ;
        RECT 116.225 135.565 116.625 135.865 ;
        RECT 115.725 134.015 116.125 134.315 ;
        RECT 115.815 133.775 116.045 134.015 ;
        RECT 116.295 133.775 116.525 135.565 ;
        RECT 116.860 134.315 117.090 141.775 ;
        RECT 117.340 136.515 117.570 141.775 ;
        RECT 117.275 136.215 117.675 136.515 ;
        RECT 116.775 134.015 117.175 134.315 ;
        RECT 116.860 133.775 117.090 134.015 ;
        RECT 117.340 133.775 117.570 136.215 ;
        RECT 117.820 134.315 118.050 141.775 ;
        RECT 118.300 136.515 118.530 141.775 ;
        RECT 118.225 136.215 118.625 136.515 ;
        RECT 117.725 134.015 118.125 134.315 ;
        RECT 117.820 133.775 118.050 134.015 ;
        RECT 118.300 133.775 118.530 136.215 ;
        RECT 118.780 134.315 119.010 141.775 ;
        RECT 119.260 136.515 119.490 141.775 ;
        RECT 119.175 136.215 119.575 136.515 ;
        RECT 118.675 134.015 119.075 134.315 ;
        RECT 118.780 133.775 119.010 134.015 ;
        RECT 119.260 133.775 119.490 136.215 ;
        RECT 119.740 134.315 119.970 141.775 ;
        RECT 120.220 136.515 120.450 141.775 ;
        RECT 120.125 136.215 120.525 136.515 ;
        RECT 119.675 134.015 120.075 134.315 ;
        RECT 119.740 133.775 119.970 134.015 ;
        RECT 120.220 133.775 120.450 136.215 ;
        RECT 120.700 134.315 120.930 141.775 ;
        RECT 121.180 136.515 121.410 141.775 ;
        RECT 121.075 136.215 121.475 136.515 ;
        RECT 120.625 134.015 121.025 134.315 ;
        RECT 120.700 133.775 120.930 134.015 ;
        RECT 121.180 133.775 121.410 136.215 ;
        RECT 121.660 134.315 121.890 141.775 ;
        RECT 122.140 136.515 122.370 141.775 ;
        RECT 122.075 136.215 122.475 136.515 ;
        RECT 121.575 134.015 121.975 134.315 ;
        RECT 121.660 133.775 121.890 134.015 ;
        RECT 122.140 133.775 122.370 136.215 ;
        RECT 122.620 134.315 122.850 141.775 ;
        RECT 123.100 136.515 123.330 141.775 ;
        RECT 123.025 136.215 123.425 136.515 ;
        RECT 122.525 134.015 122.925 134.315 ;
        RECT 122.620 133.775 122.850 134.015 ;
        RECT 123.100 133.775 123.330 136.215 ;
        RECT 123.580 134.315 123.810 141.775 ;
        RECT 124.060 136.515 124.290 141.775 ;
        RECT 123.975 136.215 124.375 136.515 ;
        RECT 123.475 134.015 123.875 134.315 ;
        RECT 123.580 133.775 123.810 134.015 ;
        RECT 124.060 133.775 124.290 136.215 ;
        RECT 124.675 133.415 125.025 142.565 ;
        RECT 85.825 133.065 125.025 133.415 ;
        RECT 125.175 142.565 153.825 142.915 ;
        RECT 125.175 133.415 125.425 142.565 ;
        RECT 126.025 142.015 126.425 142.315 ;
        RECT 127.175 142.015 127.575 142.315 ;
        RECT 128.425 142.015 128.825 142.315 ;
        RECT 129.625 142.015 130.025 142.315 ;
        RECT 130.825 142.015 131.225 142.315 ;
        RECT 132.075 142.015 132.475 142.315 ;
        RECT 133.275 142.015 133.675 142.315 ;
        RECT 134.525 142.265 134.925 142.315 ;
        RECT 137.125 142.265 137.525 142.315 ;
        RECT 142.225 142.265 142.625 142.315 ;
        RECT 152.475 142.270 152.875 142.315 ;
        RECT 133.925 142.015 134.975 142.265 ;
        RECT 135.175 142.015 137.525 142.265 ;
        RECT 137.725 142.015 142.675 142.265 ;
        RECT 142.875 142.020 152.875 142.270 ;
        RECT 152.475 142.015 152.875 142.020 ;
        RECT 125.765 137.815 125.995 141.815 ;
        RECT 126.405 138.565 126.635 141.815 ;
        RECT 126.325 138.265 126.725 138.565 ;
        RECT 126.405 137.815 126.635 138.265 ;
        RECT 126.975 137.815 127.205 141.815 ;
        RECT 127.615 138.565 127.845 141.815 ;
        RECT 127.525 138.265 127.925 138.565 ;
        RECT 128.185 138.265 128.415 141.815 ;
        RECT 128.825 138.565 129.055 141.815 ;
        RECT 128.725 138.265 129.125 138.565 ;
        RECT 127.615 137.815 127.845 138.265 ;
        RECT 128.175 137.815 128.415 138.265 ;
        RECT 128.825 137.815 129.055 138.265 ;
        RECT 129.395 137.815 129.625 141.815 ;
        RECT 130.035 138.565 130.265 141.815 ;
        RECT 129.975 138.265 130.375 138.565 ;
        RECT 130.035 137.815 130.265 138.265 ;
        RECT 130.605 137.815 130.835 141.815 ;
        RECT 131.245 138.565 131.475 141.815 ;
        RECT 131.175 138.265 131.575 138.565 ;
        RECT 131.245 137.815 131.475 138.265 ;
        RECT 131.815 137.815 132.045 141.815 ;
        RECT 132.455 138.565 132.685 141.815 ;
        RECT 132.375 138.265 132.775 138.565 ;
        RECT 132.455 137.815 132.685 138.265 ;
        RECT 125.775 134.065 125.975 137.815 ;
        RECT 126.975 134.065 127.175 137.815 ;
        RECT 128.175 134.065 128.375 137.815 ;
        RECT 129.425 134.065 129.625 137.815 ;
        RECT 130.625 134.065 130.825 137.815 ;
        RECT 131.825 134.065 132.025 137.815 ;
        RECT 133.040 134.215 133.270 141.815 ;
        RECT 133.680 138.565 133.910 141.815 ;
        RECT 133.575 138.265 133.975 138.565 ;
        RECT 125.675 133.765 126.075 134.065 ;
        RECT 126.875 133.765 127.275 134.065 ;
        RECT 128.075 133.765 128.475 134.065 ;
        RECT 129.325 133.765 129.725 134.065 ;
        RECT 130.525 133.765 130.925 134.065 ;
        RECT 131.725 133.765 132.125 134.065 ;
        RECT 132.975 133.915 133.375 134.215 ;
        RECT 133.040 133.815 133.270 133.915 ;
        RECT 133.680 133.815 133.910 138.265 ;
        RECT 134.320 134.215 134.550 141.815 ;
        RECT 134.960 138.565 135.190 141.815 ;
        RECT 134.875 138.265 135.275 138.565 ;
        RECT 134.225 133.915 134.625 134.215 ;
        RECT 134.320 133.815 134.550 133.915 ;
        RECT 134.960 133.815 135.190 138.265 ;
        RECT 135.600 134.215 135.830 141.815 ;
        RECT 136.240 138.565 136.470 141.815 ;
        RECT 136.175 138.265 136.575 138.565 ;
        RECT 135.525 133.915 135.925 134.215 ;
        RECT 135.600 133.815 135.830 133.915 ;
        RECT 136.240 133.815 136.470 138.265 ;
        RECT 136.880 134.215 137.110 141.815 ;
        RECT 137.520 138.565 137.750 141.815 ;
        RECT 137.425 138.265 137.825 138.565 ;
        RECT 136.825 133.915 137.225 134.215 ;
        RECT 136.880 133.815 137.110 133.915 ;
        RECT 137.520 133.815 137.750 138.265 ;
        RECT 138.160 134.215 138.390 141.815 ;
        RECT 138.800 138.565 139.030 141.815 ;
        RECT 138.725 138.265 139.125 138.565 ;
        RECT 138.075 133.915 138.475 134.215 ;
        RECT 138.160 133.815 138.390 133.915 ;
        RECT 138.800 133.815 139.030 138.265 ;
        RECT 139.440 134.215 139.670 141.815 ;
        RECT 140.080 138.565 140.310 141.815 ;
        RECT 140.025 138.265 140.425 138.565 ;
        RECT 139.375 133.915 139.775 134.215 ;
        RECT 139.440 133.815 139.670 133.915 ;
        RECT 140.080 133.815 140.310 138.265 ;
        RECT 140.720 134.215 140.950 141.815 ;
        RECT 141.360 138.565 141.590 141.815 ;
        RECT 141.275 138.265 141.675 138.565 ;
        RECT 140.625 133.915 141.025 134.215 ;
        RECT 140.720 133.815 140.950 133.915 ;
        RECT 141.360 133.815 141.590 138.265 ;
        RECT 142.000 134.215 142.230 141.815 ;
        RECT 142.640 138.565 142.870 141.815 ;
        RECT 142.575 138.265 142.975 138.565 ;
        RECT 141.925 133.915 142.325 134.215 ;
        RECT 142.000 133.815 142.230 133.915 ;
        RECT 142.640 133.815 142.870 138.265 ;
        RECT 143.280 134.215 143.510 141.815 ;
        RECT 143.920 138.565 144.150 141.815 ;
        RECT 143.825 138.265 144.225 138.565 ;
        RECT 143.175 133.915 143.575 134.215 ;
        RECT 143.280 133.815 143.510 133.915 ;
        RECT 143.920 133.815 144.150 138.265 ;
        RECT 144.560 134.215 144.790 141.815 ;
        RECT 145.200 138.565 145.430 141.815 ;
        RECT 145.125 138.265 145.525 138.565 ;
        RECT 144.475 133.915 144.875 134.215 ;
        RECT 144.560 133.815 144.790 133.915 ;
        RECT 145.200 133.815 145.430 138.265 ;
        RECT 145.840 134.215 146.070 141.815 ;
        RECT 146.480 138.565 146.710 141.815 ;
        RECT 146.425 138.265 146.825 138.565 ;
        RECT 145.775 133.915 146.175 134.215 ;
        RECT 145.840 133.815 146.070 133.915 ;
        RECT 146.480 133.815 146.710 138.265 ;
        RECT 147.120 134.215 147.350 141.815 ;
        RECT 147.760 138.565 147.990 141.815 ;
        RECT 147.675 138.265 148.075 138.565 ;
        RECT 147.025 133.915 147.425 134.215 ;
        RECT 147.120 133.815 147.350 133.915 ;
        RECT 147.760 133.815 147.990 138.265 ;
        RECT 148.400 134.215 148.630 141.815 ;
        RECT 149.040 138.565 149.270 141.815 ;
        RECT 148.975 138.265 149.375 138.565 ;
        RECT 148.325 133.915 148.725 134.215 ;
        RECT 148.400 133.815 148.630 133.915 ;
        RECT 149.040 133.815 149.270 138.265 ;
        RECT 149.680 134.215 149.910 141.815 ;
        RECT 150.320 138.565 150.550 141.815 ;
        RECT 150.225 138.265 150.625 138.565 ;
        RECT 149.575 133.915 149.975 134.215 ;
        RECT 149.680 133.815 149.910 133.915 ;
        RECT 150.320 133.815 150.550 138.265 ;
        RECT 150.960 134.215 151.190 141.815 ;
        RECT 151.600 138.565 151.830 141.815 ;
        RECT 151.525 138.265 151.925 138.565 ;
        RECT 150.875 133.915 151.275 134.215 ;
        RECT 150.960 133.815 151.190 133.915 ;
        RECT 151.600 133.815 151.830 138.265 ;
        RECT 152.240 134.215 152.470 141.815 ;
        RECT 152.880 138.565 153.110 141.815 ;
        RECT 152.825 138.265 153.225 138.565 ;
        RECT 152.175 133.915 152.575 134.215 ;
        RECT 152.240 133.815 152.470 133.915 ;
        RECT 152.880 133.815 153.110 138.265 ;
        RECT 153.425 133.415 153.825 142.565 ;
        RECT 125.175 133.065 153.825 133.415 ;
        RECT 8.540 132.615 8.940 132.690 ;
        RECT 37.240 132.615 37.640 132.690 ;
        RECT 44.990 132.615 45.390 132.690 ;
        RECT 50.890 132.615 51.290 132.690 ;
        RECT 74.940 132.615 75.340 132.690 ;
        RECT 8.540 132.465 75.340 132.615 ;
        RECT 8.540 132.390 8.940 132.465 ;
        RECT 37.240 132.390 37.640 132.465 ;
        RECT 44.990 132.390 45.390 132.465 ;
        RECT 50.890 132.390 51.290 132.465 ;
        RECT 74.940 132.390 75.340 132.465 ;
        RECT 85.775 132.615 86.175 132.690 ;
        RECT 109.825 132.615 110.225 132.690 ;
        RECT 115.725 132.615 116.125 132.690 ;
        RECT 123.475 132.615 123.875 132.690 ;
        RECT 152.175 132.615 152.575 132.690 ;
        RECT 85.775 132.465 152.575 132.615 ;
        RECT 85.775 132.390 86.175 132.465 ;
        RECT 109.825 132.390 110.225 132.465 ;
        RECT 115.725 132.390 116.125 132.465 ;
        RECT 123.475 132.390 123.875 132.465 ;
        RECT 152.175 132.390 152.575 132.465 ;
        RECT 18.790 132.165 19.190 132.240 ;
        RECT 41.040 132.165 41.440 132.240 ;
        RECT 45.940 132.165 46.340 132.240 ;
        RECT 54.740 132.165 55.140 132.240 ;
        RECT 75.390 132.165 75.790 132.240 ;
        RECT 18.790 132.015 75.790 132.165 ;
        RECT 18.790 131.940 19.190 132.015 ;
        RECT 41.040 131.940 41.440 132.015 ;
        RECT 45.940 131.940 46.340 132.015 ;
        RECT 54.740 131.940 55.140 132.015 ;
        RECT 75.390 131.940 75.790 132.015 ;
        RECT 85.325 132.165 85.725 132.240 ;
        RECT 105.975 132.165 106.375 132.240 ;
        RECT 114.775 132.165 115.175 132.240 ;
        RECT 119.675 132.165 120.075 132.240 ;
        RECT 141.925 132.165 142.325 132.240 ;
        RECT 85.325 132.015 142.325 132.165 ;
        RECT 85.325 131.940 85.725 132.015 ;
        RECT 105.975 131.940 106.375 132.015 ;
        RECT 114.775 131.940 115.175 132.015 ;
        RECT 119.675 131.940 120.075 132.015 ;
        RECT 141.925 131.940 142.325 132.015 ;
        RECT 23.890 131.715 24.290 131.790 ;
        RECT 42.990 131.715 43.390 131.790 ;
        RECT 56.640 131.715 57.040 131.790 ;
        RECT 66.990 131.715 67.390 131.790 ;
        RECT 75.840 131.715 76.240 131.790 ;
        RECT 23.890 131.565 76.240 131.715 ;
        RECT 23.890 131.490 24.290 131.565 ;
        RECT 42.990 131.490 43.390 131.565 ;
        RECT 56.640 131.490 57.040 131.565 ;
        RECT 66.990 131.490 67.390 131.565 ;
        RECT 75.840 131.490 76.240 131.565 ;
        RECT 84.875 131.715 85.275 131.790 ;
        RECT 93.725 131.715 94.125 131.790 ;
        RECT 104.075 131.715 104.475 131.790 ;
        RECT 117.725 131.715 118.125 131.790 ;
        RECT 136.825 131.715 137.225 131.790 ;
        RECT 84.875 131.565 137.225 131.715 ;
        RECT 84.875 131.490 85.275 131.565 ;
        RECT 93.725 131.490 94.125 131.565 ;
        RECT 104.075 131.490 104.475 131.565 ;
        RECT 117.725 131.490 118.125 131.565 ;
        RECT 136.825 131.490 137.225 131.565 ;
        RECT 26.490 131.265 26.890 131.340 ;
        RECT 43.940 131.265 44.340 131.340 ;
        RECT 57.640 131.265 58.040 131.340 ;
        RECT 67.940 131.265 68.340 131.340 ;
        RECT 76.290 131.265 76.690 131.340 ;
        RECT 26.490 131.115 76.690 131.265 ;
        RECT 26.490 131.040 26.890 131.115 ;
        RECT 43.940 131.040 44.340 131.115 ;
        RECT 57.640 131.040 58.040 131.115 ;
        RECT 67.940 131.040 68.340 131.115 ;
        RECT 76.290 131.040 76.690 131.115 ;
        RECT 84.425 131.265 84.825 131.340 ;
        RECT 92.775 131.265 93.175 131.340 ;
        RECT 103.075 131.265 103.475 131.340 ;
        RECT 116.775 131.265 117.175 131.340 ;
        RECT 134.225 131.265 134.625 131.340 ;
        RECT 84.425 131.115 134.625 131.265 ;
        RECT 84.425 131.040 84.825 131.115 ;
        RECT 92.775 131.040 93.175 131.115 ;
        RECT 103.075 131.040 103.475 131.115 ;
        RECT 116.775 131.040 117.175 131.115 ;
        RECT 134.225 131.040 134.625 131.115 ;
        RECT 27.740 130.815 28.140 130.890 ;
        RECT 58.690 130.815 59.090 130.890 ;
        RECT 68.490 130.815 68.890 130.890 ;
        RECT 76.740 130.815 77.140 130.890 ;
        RECT 27.740 130.665 77.140 130.815 ;
        RECT 27.740 130.590 28.140 130.665 ;
        RECT 58.690 130.590 59.090 130.665 ;
        RECT 68.490 130.590 68.890 130.665 ;
        RECT 76.740 130.590 77.140 130.665 ;
        RECT 83.975 130.815 84.375 130.890 ;
        RECT 92.225 130.815 92.625 130.890 ;
        RECT 102.025 130.815 102.425 130.890 ;
        RECT 132.975 130.815 133.375 130.890 ;
        RECT 83.975 130.665 133.375 130.815 ;
        RECT 83.975 130.590 84.375 130.665 ;
        RECT 92.225 130.590 92.625 130.665 ;
        RECT 102.025 130.590 102.425 130.665 ;
        RECT 132.975 130.590 133.375 130.665 ;
        RECT 28.990 130.365 29.390 130.440 ;
        RECT 59.640 130.365 60.040 130.440 ;
        RECT 69.540 130.365 69.940 130.440 ;
        RECT 77.190 130.365 77.590 130.440 ;
        RECT 28.990 130.215 77.590 130.365 ;
        RECT 28.990 130.140 29.390 130.215 ;
        RECT 59.640 130.140 60.040 130.215 ;
        RECT 69.540 130.140 69.940 130.215 ;
        RECT 77.190 130.140 77.590 130.215 ;
        RECT 83.525 130.365 83.925 130.440 ;
        RECT 91.175 130.365 91.575 130.440 ;
        RECT 101.075 130.365 101.475 130.440 ;
        RECT 131.725 130.365 132.125 130.440 ;
        RECT 83.525 130.215 132.125 130.365 ;
        RECT 83.525 130.140 83.925 130.215 ;
        RECT 91.175 130.140 91.575 130.215 ;
        RECT 101.075 130.140 101.475 130.215 ;
        RECT 131.725 130.140 132.125 130.215 ;
        RECT 30.190 129.915 30.590 129.990 ;
        RECT 60.690 129.915 61.090 129.990 ;
        RECT 70.590 129.915 70.990 129.990 ;
        RECT 77.640 129.915 78.040 129.990 ;
        RECT 30.190 129.765 78.040 129.915 ;
        RECT 30.190 129.690 30.590 129.765 ;
        RECT 60.690 129.690 61.090 129.765 ;
        RECT 70.590 129.690 70.990 129.765 ;
        RECT 77.640 129.690 78.040 129.765 ;
        RECT 83.075 129.915 83.475 129.990 ;
        RECT 90.125 129.915 90.525 129.990 ;
        RECT 100.025 129.915 100.425 129.990 ;
        RECT 130.525 129.915 130.925 129.990 ;
        RECT 83.075 129.765 130.925 129.915 ;
        RECT 83.075 129.690 83.475 129.765 ;
        RECT 90.125 129.690 90.525 129.765 ;
        RECT 100.025 129.690 100.425 129.765 ;
        RECT 130.525 129.690 130.925 129.765 ;
        RECT 31.390 129.465 31.790 129.540 ;
        RECT 61.740 129.465 62.140 129.540 ;
        RECT 73.640 129.465 74.040 129.540 ;
        RECT 79.890 129.465 80.290 129.540 ;
        RECT 31.390 129.315 80.290 129.465 ;
        RECT 31.390 129.240 31.790 129.315 ;
        RECT 61.740 129.240 62.140 129.315 ;
        RECT 73.640 129.240 74.040 129.315 ;
        RECT 79.890 129.240 80.290 129.315 ;
        RECT 80.825 129.465 81.225 129.540 ;
        RECT 87.075 129.465 87.475 129.540 ;
        RECT 98.975 129.465 99.375 129.540 ;
        RECT 129.325 129.465 129.725 129.540 ;
        RECT 80.825 129.315 129.725 129.465 ;
        RECT 80.825 129.240 81.225 129.315 ;
        RECT 87.075 129.240 87.475 129.315 ;
        RECT 98.975 129.240 99.375 129.315 ;
        RECT 129.325 129.240 129.725 129.315 ;
        RECT 32.640 129.015 33.040 129.090 ;
        RECT 62.790 129.015 63.190 129.090 ;
        RECT 71.640 129.015 72.040 129.090 ;
        RECT 78.090 129.015 78.490 129.090 ;
        RECT 32.640 128.865 78.490 129.015 ;
        RECT 32.640 128.790 33.040 128.865 ;
        RECT 62.790 128.790 63.190 128.865 ;
        RECT 71.640 128.790 72.040 128.865 ;
        RECT 78.090 128.790 78.490 128.865 ;
        RECT 82.625 129.015 83.025 129.090 ;
        RECT 89.075 129.015 89.475 129.090 ;
        RECT 97.925 129.015 98.325 129.090 ;
        RECT 128.075 129.015 128.475 129.090 ;
        RECT 82.625 128.865 128.475 129.015 ;
        RECT 82.625 128.790 83.025 128.865 ;
        RECT 89.075 128.790 89.475 128.865 ;
        RECT 97.925 128.790 98.325 128.865 ;
        RECT 128.075 128.790 128.475 128.865 ;
        RECT 33.840 128.565 34.240 128.640 ;
        RECT 63.840 128.565 64.240 128.640 ;
        RECT 74.040 128.565 74.440 128.640 ;
        RECT 79.440 128.565 79.840 128.640 ;
        RECT 33.840 128.415 79.840 128.565 ;
        RECT 33.840 128.340 34.240 128.415 ;
        RECT 63.840 128.340 64.240 128.415 ;
        RECT 74.040 128.340 74.440 128.415 ;
        RECT 79.440 128.340 79.840 128.415 ;
        RECT 81.275 128.565 81.675 128.640 ;
        RECT 86.675 128.565 87.075 128.640 ;
        RECT 96.875 128.565 97.275 128.640 ;
        RECT 126.875 128.565 127.275 128.640 ;
        RECT 81.275 128.415 127.275 128.565 ;
        RECT 81.275 128.340 81.675 128.415 ;
        RECT 86.675 128.340 87.075 128.415 ;
        RECT 96.875 128.340 97.275 128.415 ;
        RECT 126.875 128.340 127.275 128.415 ;
        RECT 35.040 128.115 35.440 128.190 ;
        RECT 64.890 128.115 65.290 128.190 ;
        RECT 72.690 128.115 73.090 128.190 ;
        RECT 78.990 128.115 79.390 128.190 ;
        RECT 35.040 127.965 79.390 128.115 ;
        RECT 35.040 127.890 35.440 127.965 ;
        RECT 64.890 127.890 65.290 127.965 ;
        RECT 72.690 127.890 73.090 127.965 ;
        RECT 78.990 127.890 79.390 127.965 ;
        RECT 81.725 128.115 82.125 128.190 ;
        RECT 88.025 128.115 88.425 128.190 ;
        RECT 95.825 128.115 96.225 128.190 ;
        RECT 125.675 128.115 126.075 128.190 ;
        RECT 81.725 127.965 126.075 128.115 ;
        RECT 81.725 127.890 82.125 127.965 ;
        RECT 88.025 127.890 88.425 127.965 ;
        RECT 95.825 127.890 96.225 127.965 ;
        RECT 125.675 127.890 126.075 127.965 ;
        RECT 65.940 127.665 66.340 127.740 ;
        RECT 74.440 127.665 74.840 127.740 ;
        RECT 78.540 127.665 78.940 127.740 ;
        RECT 7.390 127.240 8.290 127.540 ;
        RECT 65.940 127.515 78.940 127.665 ;
        RECT 65.940 127.440 66.340 127.515 ;
        RECT 74.440 127.440 74.840 127.515 ;
        RECT 78.540 127.440 78.940 127.515 ;
        RECT 82.175 127.665 82.575 127.740 ;
        RECT 86.275 127.665 86.675 127.740 ;
        RECT 94.775 127.665 95.175 127.740 ;
        RECT 82.175 127.515 95.175 127.665 ;
        RECT 82.175 127.440 82.575 127.515 ;
        RECT 86.275 127.440 86.675 127.515 ;
        RECT 94.775 127.440 95.175 127.515 ;
        RECT 6.890 126.040 7.290 126.440 ;
        RECT 7.740 126.070 7.940 127.240 ;
        RECT 73.390 126.990 74.290 127.290 ;
        RECT 86.825 126.990 87.725 127.290 ;
        RECT 152.825 127.240 153.725 127.540 ;
        RECT 8.890 126.070 9.290 126.440 ;
        RECT 10.890 126.070 11.290 126.440 ;
        RECT 12.890 126.070 13.290 126.440 ;
        RECT 14.890 126.070 15.290 126.440 ;
        RECT 16.890 126.070 17.290 126.440 ;
        RECT 18.890 126.070 19.290 126.440 ;
        RECT 20.890 126.070 21.290 126.440 ;
        RECT 22.890 126.070 23.290 126.440 ;
        RECT 24.890 126.070 25.290 126.440 ;
        RECT 26.890 126.070 27.290 126.440 ;
        RECT 28.890 126.070 29.290 126.440 ;
        RECT 30.890 126.070 31.290 126.440 ;
        RECT 32.890 126.070 33.290 126.440 ;
        RECT 34.890 126.070 35.290 126.440 ;
        RECT 36.890 126.070 37.290 126.440 ;
        RECT 38.890 126.070 39.290 126.440 ;
        RECT 40.890 126.070 41.290 126.440 ;
        RECT 42.890 126.070 43.290 126.440 ;
        RECT 44.890 126.070 45.290 126.440 ;
        RECT 46.890 126.070 47.290 126.440 ;
        RECT 48.890 126.070 49.290 126.440 ;
        RECT 50.890 126.070 51.290 126.440 ;
        RECT 52.890 126.070 53.290 126.440 ;
        RECT 54.890 126.070 55.290 126.440 ;
        RECT 56.890 126.070 57.290 126.440 ;
        RECT 58.890 126.070 59.290 126.440 ;
        RECT 60.890 126.070 61.290 126.440 ;
        RECT 62.890 126.070 63.290 126.440 ;
        RECT 64.890 126.070 65.290 126.440 ;
        RECT 66.890 126.070 67.290 126.440 ;
        RECT 68.890 126.070 69.290 126.440 ;
        RECT 70.890 126.070 71.290 126.440 ;
        RECT 72.890 126.070 73.290 126.440 ;
        RECT 7.430 126.040 73.450 126.070 ;
        RECT 73.740 126.040 73.940 126.990 ;
        RECT 87.175 126.040 87.375 126.990 ;
        RECT 87.825 126.070 88.225 126.440 ;
        RECT 89.825 126.070 90.225 126.440 ;
        RECT 91.825 126.070 92.225 126.440 ;
        RECT 93.825 126.070 94.225 126.440 ;
        RECT 95.825 126.070 96.225 126.440 ;
        RECT 97.825 126.070 98.225 126.440 ;
        RECT 99.825 126.070 100.225 126.440 ;
        RECT 101.825 126.070 102.225 126.440 ;
        RECT 103.825 126.070 104.225 126.440 ;
        RECT 105.825 126.070 106.225 126.440 ;
        RECT 107.825 126.070 108.225 126.440 ;
        RECT 109.825 126.070 110.225 126.440 ;
        RECT 111.825 126.070 112.225 126.440 ;
        RECT 113.825 126.070 114.225 126.440 ;
        RECT 115.825 126.070 116.225 126.440 ;
        RECT 117.825 126.070 118.225 126.440 ;
        RECT 119.825 126.070 120.225 126.440 ;
        RECT 121.825 126.070 122.225 126.440 ;
        RECT 123.825 126.070 124.225 126.440 ;
        RECT 125.825 126.070 126.225 126.440 ;
        RECT 127.825 126.070 128.225 126.440 ;
        RECT 129.825 126.070 130.225 126.440 ;
        RECT 131.825 126.070 132.225 126.440 ;
        RECT 133.825 126.070 134.225 126.440 ;
        RECT 135.825 126.070 136.225 126.440 ;
        RECT 137.825 126.070 138.225 126.440 ;
        RECT 139.825 126.070 140.225 126.440 ;
        RECT 141.825 126.070 142.225 126.440 ;
        RECT 143.825 126.070 144.225 126.440 ;
        RECT 145.825 126.070 146.225 126.440 ;
        RECT 147.825 126.070 148.225 126.440 ;
        RECT 149.825 126.070 150.225 126.440 ;
        RECT 151.825 126.070 152.225 126.440 ;
        RECT 153.175 126.070 153.375 127.240 ;
        RECT 87.665 126.040 153.685 126.070 ;
        RECT 153.825 126.040 154.225 126.440 ;
        RECT 6.890 125.840 74.540 126.040 ;
        RECT 86.575 125.840 154.225 126.040 ;
        RECT 6.890 125.440 7.290 125.840 ;
        RECT 7.430 125.810 73.450 125.840 ;
        RECT 87.665 125.810 153.685 125.840 ;
        RECT 8.890 125.440 9.290 125.810 ;
        RECT 10.890 125.440 11.290 125.810 ;
        RECT 12.890 125.440 13.290 125.810 ;
        RECT 14.890 125.440 15.290 125.810 ;
        RECT 16.890 125.440 17.290 125.810 ;
        RECT 18.890 125.440 19.290 125.810 ;
        RECT 20.890 125.440 21.290 125.810 ;
        RECT 22.890 125.440 23.290 125.810 ;
        RECT 24.890 125.440 25.290 125.810 ;
        RECT 26.890 125.440 27.290 125.810 ;
        RECT 28.890 125.440 29.290 125.810 ;
        RECT 30.890 125.440 31.290 125.810 ;
        RECT 32.890 125.440 33.290 125.810 ;
        RECT 34.890 125.440 35.290 125.810 ;
        RECT 36.890 125.440 37.290 125.810 ;
        RECT 38.890 125.440 39.290 125.810 ;
        RECT 40.890 125.440 41.290 125.810 ;
        RECT 42.890 125.440 43.290 125.810 ;
        RECT 44.890 125.440 45.290 125.810 ;
        RECT 46.890 125.440 47.290 125.810 ;
        RECT 48.890 125.440 49.290 125.810 ;
        RECT 50.890 125.440 51.290 125.810 ;
        RECT 52.890 125.440 53.290 125.810 ;
        RECT 54.890 125.440 55.290 125.810 ;
        RECT 56.890 125.440 57.290 125.810 ;
        RECT 58.890 125.440 59.290 125.810 ;
        RECT 60.890 125.440 61.290 125.810 ;
        RECT 62.890 125.440 63.290 125.810 ;
        RECT 64.890 125.440 65.290 125.810 ;
        RECT 66.890 125.440 67.290 125.810 ;
        RECT 68.890 125.440 69.290 125.810 ;
        RECT 70.890 125.440 71.290 125.810 ;
        RECT 72.890 125.440 73.290 125.810 ;
        RECT 87.825 125.440 88.225 125.810 ;
        RECT 89.825 125.440 90.225 125.810 ;
        RECT 91.825 125.440 92.225 125.810 ;
        RECT 93.825 125.440 94.225 125.810 ;
        RECT 95.825 125.440 96.225 125.810 ;
        RECT 97.825 125.440 98.225 125.810 ;
        RECT 99.825 125.440 100.225 125.810 ;
        RECT 101.825 125.440 102.225 125.810 ;
        RECT 103.825 125.440 104.225 125.810 ;
        RECT 105.825 125.440 106.225 125.810 ;
        RECT 107.825 125.440 108.225 125.810 ;
        RECT 109.825 125.440 110.225 125.810 ;
        RECT 111.825 125.440 112.225 125.810 ;
        RECT 113.825 125.440 114.225 125.810 ;
        RECT 115.825 125.440 116.225 125.810 ;
        RECT 117.825 125.440 118.225 125.810 ;
        RECT 119.825 125.440 120.225 125.810 ;
        RECT 121.825 125.440 122.225 125.810 ;
        RECT 123.825 125.440 124.225 125.810 ;
        RECT 125.825 125.440 126.225 125.810 ;
        RECT 127.825 125.440 128.225 125.810 ;
        RECT 129.825 125.440 130.225 125.810 ;
        RECT 131.825 125.440 132.225 125.810 ;
        RECT 133.825 125.440 134.225 125.810 ;
        RECT 135.825 125.440 136.225 125.810 ;
        RECT 137.825 125.440 138.225 125.810 ;
        RECT 139.825 125.440 140.225 125.810 ;
        RECT 141.825 125.440 142.225 125.810 ;
        RECT 143.825 125.440 144.225 125.810 ;
        RECT 145.825 125.440 146.225 125.810 ;
        RECT 147.825 125.440 148.225 125.810 ;
        RECT 149.825 125.440 150.225 125.810 ;
        RECT 151.825 125.440 152.225 125.810 ;
        RECT 153.825 125.440 154.225 125.840 ;
        RECT 6.960 124.590 7.220 125.440 ;
        RECT 153.895 124.590 154.155 125.440 ;
        RECT 6.890 124.190 7.290 124.590 ;
        RECT 8.890 124.190 9.290 124.590 ;
        RECT 10.890 124.190 11.290 124.590 ;
        RECT 12.890 124.190 13.290 124.590 ;
        RECT 14.890 124.190 15.290 124.590 ;
        RECT 16.890 124.190 17.290 124.590 ;
        RECT 18.890 124.190 19.290 124.590 ;
        RECT 20.890 124.190 21.290 124.590 ;
        RECT 22.890 124.190 23.290 124.590 ;
        RECT 24.890 124.190 25.290 124.590 ;
        RECT 26.890 124.190 27.290 124.590 ;
        RECT 28.890 124.190 29.290 124.590 ;
        RECT 30.890 124.190 31.290 124.590 ;
        RECT 32.890 124.190 33.290 124.590 ;
        RECT 34.890 124.190 35.290 124.590 ;
        RECT 36.890 124.190 37.290 124.590 ;
        RECT 38.890 124.190 39.290 124.590 ;
        RECT 40.890 124.190 41.290 124.590 ;
        RECT 42.890 124.190 43.290 124.590 ;
        RECT 44.890 124.190 45.290 124.590 ;
        RECT 46.890 124.190 47.290 124.590 ;
        RECT 48.890 124.190 49.290 124.590 ;
        RECT 50.890 124.190 51.290 124.590 ;
        RECT 52.890 124.190 53.290 124.590 ;
        RECT 54.890 124.190 55.290 124.590 ;
        RECT 56.890 124.190 57.290 124.590 ;
        RECT 58.890 124.190 59.290 124.590 ;
        RECT 60.890 124.190 61.290 124.590 ;
        RECT 62.890 124.190 63.290 124.590 ;
        RECT 64.890 124.190 65.290 124.590 ;
        RECT 66.890 124.190 67.290 124.590 ;
        RECT 68.890 124.190 69.290 124.590 ;
        RECT 70.890 124.190 71.290 124.590 ;
        RECT 72.890 124.190 73.290 124.590 ;
        RECT 87.825 124.190 88.225 124.590 ;
        RECT 89.825 124.190 90.225 124.590 ;
        RECT 91.825 124.190 92.225 124.590 ;
        RECT 93.825 124.190 94.225 124.590 ;
        RECT 95.825 124.190 96.225 124.590 ;
        RECT 97.825 124.190 98.225 124.590 ;
        RECT 99.825 124.190 100.225 124.590 ;
        RECT 101.825 124.190 102.225 124.590 ;
        RECT 103.825 124.190 104.225 124.590 ;
        RECT 105.825 124.190 106.225 124.590 ;
        RECT 107.825 124.190 108.225 124.590 ;
        RECT 109.825 124.190 110.225 124.590 ;
        RECT 111.825 124.190 112.225 124.590 ;
        RECT 113.825 124.190 114.225 124.590 ;
        RECT 115.825 124.190 116.225 124.590 ;
        RECT 117.825 124.190 118.225 124.590 ;
        RECT 119.825 124.190 120.225 124.590 ;
        RECT 121.825 124.190 122.225 124.590 ;
        RECT 123.825 124.190 124.225 124.590 ;
        RECT 125.825 124.190 126.225 124.590 ;
        RECT 127.825 124.190 128.225 124.590 ;
        RECT 129.825 124.190 130.225 124.590 ;
        RECT 131.825 124.190 132.225 124.590 ;
        RECT 133.825 124.190 134.225 124.590 ;
        RECT 135.825 124.190 136.225 124.590 ;
        RECT 137.825 124.190 138.225 124.590 ;
        RECT 139.825 124.190 140.225 124.590 ;
        RECT 141.825 124.190 142.225 124.590 ;
        RECT 143.825 124.190 144.225 124.590 ;
        RECT 145.825 124.190 146.225 124.590 ;
        RECT 147.825 124.190 148.225 124.590 ;
        RECT 149.825 124.190 150.225 124.590 ;
        RECT 151.825 124.190 152.225 124.590 ;
        RECT 153.825 124.190 154.225 124.590 ;
        RECT 6.890 123.990 8.540 124.190 ;
        RECT 8.890 123.990 74.540 124.190 ;
        RECT 86.575 123.990 152.225 124.190 ;
        RECT 152.575 123.990 154.225 124.190 ;
        RECT 6.890 123.590 7.290 123.990 ;
        RECT 8.890 123.590 9.290 123.990 ;
        RECT 10.890 123.590 11.290 123.990 ;
        RECT 12.890 123.590 13.290 123.990 ;
        RECT 14.890 123.590 15.290 123.990 ;
        RECT 16.890 123.590 17.290 123.990 ;
        RECT 18.890 123.590 19.290 123.990 ;
        RECT 20.890 123.590 21.290 123.990 ;
        RECT 22.890 123.590 23.290 123.990 ;
        RECT 24.890 123.590 25.290 123.990 ;
        RECT 26.890 123.590 27.290 123.990 ;
        RECT 28.890 123.590 29.290 123.990 ;
        RECT 30.890 123.590 31.290 123.990 ;
        RECT 32.890 123.590 33.290 123.990 ;
        RECT 34.890 123.590 35.290 123.990 ;
        RECT 36.890 123.590 37.290 123.990 ;
        RECT 38.890 123.590 39.290 123.990 ;
        RECT 40.890 123.590 41.290 123.990 ;
        RECT 42.890 123.590 43.290 123.990 ;
        RECT 44.890 123.590 45.290 123.990 ;
        RECT 46.890 123.590 47.290 123.990 ;
        RECT 48.890 123.590 49.290 123.990 ;
        RECT 50.890 123.590 51.290 123.990 ;
        RECT 52.890 123.590 53.290 123.990 ;
        RECT 54.890 123.590 55.290 123.990 ;
        RECT 56.890 123.590 57.290 123.990 ;
        RECT 58.890 123.590 59.290 123.990 ;
        RECT 60.890 123.590 61.290 123.990 ;
        RECT 62.890 123.590 63.290 123.990 ;
        RECT 64.890 123.590 65.290 123.990 ;
        RECT 66.890 123.590 67.290 123.990 ;
        RECT 68.890 123.590 69.290 123.990 ;
        RECT 70.890 123.590 71.290 123.990 ;
        RECT 72.890 123.590 73.290 123.990 ;
        RECT 87.825 123.590 88.225 123.990 ;
        RECT 89.825 123.590 90.225 123.990 ;
        RECT 91.825 123.590 92.225 123.990 ;
        RECT 93.825 123.590 94.225 123.990 ;
        RECT 95.825 123.590 96.225 123.990 ;
        RECT 97.825 123.590 98.225 123.990 ;
        RECT 99.825 123.590 100.225 123.990 ;
        RECT 101.825 123.590 102.225 123.990 ;
        RECT 103.825 123.590 104.225 123.990 ;
        RECT 105.825 123.590 106.225 123.990 ;
        RECT 107.825 123.590 108.225 123.990 ;
        RECT 109.825 123.590 110.225 123.990 ;
        RECT 111.825 123.590 112.225 123.990 ;
        RECT 113.825 123.590 114.225 123.990 ;
        RECT 115.825 123.590 116.225 123.990 ;
        RECT 117.825 123.590 118.225 123.990 ;
        RECT 119.825 123.590 120.225 123.990 ;
        RECT 121.825 123.590 122.225 123.990 ;
        RECT 123.825 123.590 124.225 123.990 ;
        RECT 125.825 123.590 126.225 123.990 ;
        RECT 127.825 123.590 128.225 123.990 ;
        RECT 129.825 123.590 130.225 123.990 ;
        RECT 131.825 123.590 132.225 123.990 ;
        RECT 133.825 123.590 134.225 123.990 ;
        RECT 135.825 123.590 136.225 123.990 ;
        RECT 137.825 123.590 138.225 123.990 ;
        RECT 139.825 123.590 140.225 123.990 ;
        RECT 141.825 123.590 142.225 123.990 ;
        RECT 143.825 123.590 144.225 123.990 ;
        RECT 145.825 123.590 146.225 123.990 ;
        RECT 147.825 123.590 148.225 123.990 ;
        RECT 149.825 123.590 150.225 123.990 ;
        RECT 151.825 123.590 152.225 123.990 ;
        RECT 153.825 123.590 154.225 123.990 ;
        RECT 6.960 122.740 7.220 123.590 ;
        RECT 8.990 122.740 9.190 123.590 ;
        RECT 10.990 122.740 11.190 123.590 ;
        RECT 12.990 122.740 13.190 123.590 ;
        RECT 14.990 122.740 15.190 123.590 ;
        RECT 16.990 122.740 17.190 123.590 ;
        RECT 18.990 122.740 19.190 123.590 ;
        RECT 20.990 122.740 21.190 123.590 ;
        RECT 22.990 122.740 23.190 123.590 ;
        RECT 24.990 122.740 25.190 123.590 ;
        RECT 26.990 122.740 27.190 123.590 ;
        RECT 28.990 122.740 29.190 123.590 ;
        RECT 30.990 122.740 31.190 123.590 ;
        RECT 32.990 122.740 33.190 123.590 ;
        RECT 34.990 122.740 35.190 123.590 ;
        RECT 36.990 122.740 37.190 123.590 ;
        RECT 38.990 122.740 39.190 123.590 ;
        RECT 40.990 122.740 41.190 123.590 ;
        RECT 42.990 122.740 43.190 123.590 ;
        RECT 44.990 122.740 45.190 123.590 ;
        RECT 46.990 122.740 47.190 123.590 ;
        RECT 48.990 122.740 49.190 123.590 ;
        RECT 50.990 122.740 51.190 123.590 ;
        RECT 52.990 122.740 53.190 123.590 ;
        RECT 54.990 122.740 55.190 123.590 ;
        RECT 56.990 122.740 57.190 123.590 ;
        RECT 58.990 122.740 59.190 123.590 ;
        RECT 60.990 122.740 61.190 123.590 ;
        RECT 62.990 122.740 63.190 123.590 ;
        RECT 64.990 122.740 65.190 123.590 ;
        RECT 66.990 122.740 67.190 123.590 ;
        RECT 68.990 122.740 69.190 123.590 ;
        RECT 70.990 122.740 71.190 123.590 ;
        RECT 89.925 122.740 90.125 123.590 ;
        RECT 91.925 122.740 92.125 123.590 ;
        RECT 93.925 122.740 94.125 123.590 ;
        RECT 95.925 122.740 96.125 123.590 ;
        RECT 97.925 122.740 98.125 123.590 ;
        RECT 99.925 122.740 100.125 123.590 ;
        RECT 101.925 122.740 102.125 123.590 ;
        RECT 103.925 122.740 104.125 123.590 ;
        RECT 105.925 122.740 106.125 123.590 ;
        RECT 107.925 122.740 108.125 123.590 ;
        RECT 109.925 122.740 110.125 123.590 ;
        RECT 111.925 122.740 112.125 123.590 ;
        RECT 113.925 122.740 114.125 123.590 ;
        RECT 115.925 122.740 116.125 123.590 ;
        RECT 117.925 122.740 118.125 123.590 ;
        RECT 119.925 122.740 120.125 123.590 ;
        RECT 121.925 122.740 122.125 123.590 ;
        RECT 123.925 122.740 124.125 123.590 ;
        RECT 125.925 122.740 126.125 123.590 ;
        RECT 127.925 122.740 128.125 123.590 ;
        RECT 129.925 122.740 130.125 123.590 ;
        RECT 131.925 122.740 132.125 123.590 ;
        RECT 133.925 122.740 134.125 123.590 ;
        RECT 135.925 122.740 136.125 123.590 ;
        RECT 137.925 122.740 138.125 123.590 ;
        RECT 139.925 122.740 140.125 123.590 ;
        RECT 141.925 122.740 142.125 123.590 ;
        RECT 143.925 122.740 144.125 123.590 ;
        RECT 145.925 122.740 146.125 123.590 ;
        RECT 147.925 122.740 148.125 123.590 ;
        RECT 149.925 122.740 150.125 123.590 ;
        RECT 151.925 122.740 152.125 123.590 ;
        RECT 153.895 122.740 154.155 123.590 ;
        RECT 6.890 122.340 7.290 122.740 ;
        RECT 8.890 122.340 9.290 122.740 ;
        RECT 10.890 122.340 11.290 122.740 ;
        RECT 12.890 122.340 13.290 122.740 ;
        RECT 14.890 122.340 15.290 122.740 ;
        RECT 16.890 122.340 17.290 122.740 ;
        RECT 18.890 122.340 19.290 122.740 ;
        RECT 20.890 122.340 21.290 122.740 ;
        RECT 22.890 122.340 23.290 122.740 ;
        RECT 24.890 122.340 25.290 122.740 ;
        RECT 26.890 122.340 27.290 122.740 ;
        RECT 28.890 122.340 29.290 122.740 ;
        RECT 30.890 122.340 31.290 122.740 ;
        RECT 32.890 122.340 33.290 122.740 ;
        RECT 34.890 122.340 35.290 122.740 ;
        RECT 36.890 122.340 37.290 122.740 ;
        RECT 38.890 122.340 39.290 122.740 ;
        RECT 40.890 122.340 41.290 122.740 ;
        RECT 42.890 122.340 43.290 122.740 ;
        RECT 44.890 122.340 45.290 122.740 ;
        RECT 46.890 122.340 47.290 122.740 ;
        RECT 48.890 122.340 49.290 122.740 ;
        RECT 50.890 122.340 51.290 122.740 ;
        RECT 52.890 122.340 53.290 122.740 ;
        RECT 54.890 122.340 55.290 122.740 ;
        RECT 56.890 122.340 57.290 122.740 ;
        RECT 58.890 122.340 59.290 122.740 ;
        RECT 60.890 122.340 61.290 122.740 ;
        RECT 62.890 122.340 63.290 122.740 ;
        RECT 64.890 122.340 65.290 122.740 ;
        RECT 66.890 122.340 67.290 122.740 ;
        RECT 68.890 122.340 69.290 122.740 ;
        RECT 70.890 122.340 71.290 122.740 ;
        RECT 72.890 122.340 73.290 122.740 ;
        RECT 87.825 122.340 88.225 122.740 ;
        RECT 89.825 122.340 90.225 122.740 ;
        RECT 91.825 122.340 92.225 122.740 ;
        RECT 93.825 122.340 94.225 122.740 ;
        RECT 95.825 122.340 96.225 122.740 ;
        RECT 97.825 122.340 98.225 122.740 ;
        RECT 99.825 122.340 100.225 122.740 ;
        RECT 101.825 122.340 102.225 122.740 ;
        RECT 103.825 122.340 104.225 122.740 ;
        RECT 105.825 122.340 106.225 122.740 ;
        RECT 107.825 122.340 108.225 122.740 ;
        RECT 109.825 122.340 110.225 122.740 ;
        RECT 111.825 122.340 112.225 122.740 ;
        RECT 113.825 122.340 114.225 122.740 ;
        RECT 115.825 122.340 116.225 122.740 ;
        RECT 117.825 122.340 118.225 122.740 ;
        RECT 119.825 122.340 120.225 122.740 ;
        RECT 121.825 122.340 122.225 122.740 ;
        RECT 123.825 122.340 124.225 122.740 ;
        RECT 125.825 122.340 126.225 122.740 ;
        RECT 127.825 122.340 128.225 122.740 ;
        RECT 129.825 122.340 130.225 122.740 ;
        RECT 131.825 122.340 132.225 122.740 ;
        RECT 133.825 122.340 134.225 122.740 ;
        RECT 135.825 122.340 136.225 122.740 ;
        RECT 137.825 122.340 138.225 122.740 ;
        RECT 139.825 122.340 140.225 122.740 ;
        RECT 141.825 122.340 142.225 122.740 ;
        RECT 143.825 122.340 144.225 122.740 ;
        RECT 145.825 122.340 146.225 122.740 ;
        RECT 147.825 122.340 148.225 122.740 ;
        RECT 149.825 122.340 150.225 122.740 ;
        RECT 151.825 122.340 152.225 122.740 ;
        RECT 153.825 122.340 154.225 122.740 ;
        RECT 6.890 122.140 8.540 122.340 ;
        RECT 8.890 122.140 74.540 122.340 ;
        RECT 86.575 122.140 152.225 122.340 ;
        RECT 152.575 122.140 154.225 122.340 ;
        RECT 6.890 121.740 7.290 122.140 ;
        RECT 8.890 121.740 9.290 122.140 ;
        RECT 10.890 121.740 11.290 122.140 ;
        RECT 12.890 121.740 13.290 122.140 ;
        RECT 14.890 121.740 15.290 122.140 ;
        RECT 16.890 121.740 17.290 122.140 ;
        RECT 18.890 121.740 19.290 122.140 ;
        RECT 20.890 121.740 21.290 122.140 ;
        RECT 22.890 121.740 23.290 122.140 ;
        RECT 24.890 121.740 25.290 122.140 ;
        RECT 26.890 121.740 27.290 122.140 ;
        RECT 28.890 121.740 29.290 122.140 ;
        RECT 30.890 121.740 31.290 122.140 ;
        RECT 32.890 121.740 33.290 122.140 ;
        RECT 34.890 121.740 35.290 122.140 ;
        RECT 36.890 121.740 37.290 122.140 ;
        RECT 38.890 121.740 39.290 122.140 ;
        RECT 40.890 121.740 41.290 122.140 ;
        RECT 42.890 121.740 43.290 122.140 ;
        RECT 44.890 121.740 45.290 122.140 ;
        RECT 46.890 121.740 47.290 122.140 ;
        RECT 48.890 121.740 49.290 122.140 ;
        RECT 50.890 121.740 51.290 122.140 ;
        RECT 52.890 121.740 53.290 122.140 ;
        RECT 54.890 121.740 55.290 122.140 ;
        RECT 56.890 121.740 57.290 122.140 ;
        RECT 58.890 121.740 59.290 122.140 ;
        RECT 60.890 121.740 61.290 122.140 ;
        RECT 62.890 121.740 63.290 122.140 ;
        RECT 64.890 121.740 65.290 122.140 ;
        RECT 66.890 121.740 67.290 122.140 ;
        RECT 68.890 121.740 69.290 122.140 ;
        RECT 70.890 121.740 71.290 122.140 ;
        RECT 72.890 121.740 73.290 122.140 ;
        RECT 87.825 121.740 88.225 122.140 ;
        RECT 89.825 121.740 90.225 122.140 ;
        RECT 91.825 121.740 92.225 122.140 ;
        RECT 93.825 121.740 94.225 122.140 ;
        RECT 95.825 121.740 96.225 122.140 ;
        RECT 97.825 121.740 98.225 122.140 ;
        RECT 99.825 121.740 100.225 122.140 ;
        RECT 101.825 121.740 102.225 122.140 ;
        RECT 103.825 121.740 104.225 122.140 ;
        RECT 105.825 121.740 106.225 122.140 ;
        RECT 107.825 121.740 108.225 122.140 ;
        RECT 109.825 121.740 110.225 122.140 ;
        RECT 111.825 121.740 112.225 122.140 ;
        RECT 113.825 121.740 114.225 122.140 ;
        RECT 115.825 121.740 116.225 122.140 ;
        RECT 117.825 121.740 118.225 122.140 ;
        RECT 119.825 121.740 120.225 122.140 ;
        RECT 121.825 121.740 122.225 122.140 ;
        RECT 123.825 121.740 124.225 122.140 ;
        RECT 125.825 121.740 126.225 122.140 ;
        RECT 127.825 121.740 128.225 122.140 ;
        RECT 129.825 121.740 130.225 122.140 ;
        RECT 131.825 121.740 132.225 122.140 ;
        RECT 133.825 121.740 134.225 122.140 ;
        RECT 135.825 121.740 136.225 122.140 ;
        RECT 137.825 121.740 138.225 122.140 ;
        RECT 139.825 121.740 140.225 122.140 ;
        RECT 141.825 121.740 142.225 122.140 ;
        RECT 143.825 121.740 144.225 122.140 ;
        RECT 145.825 121.740 146.225 122.140 ;
        RECT 147.825 121.740 148.225 122.140 ;
        RECT 149.825 121.740 150.225 122.140 ;
        RECT 151.825 121.740 152.225 122.140 ;
        RECT 153.825 121.740 154.225 122.140 ;
        RECT 6.960 120.890 7.220 121.740 ;
        RECT 8.990 120.890 9.190 121.740 ;
        RECT 10.990 120.890 11.190 121.740 ;
        RECT 12.990 120.890 13.190 121.740 ;
        RECT 14.990 120.890 15.190 121.740 ;
        RECT 16.990 120.890 17.190 121.740 ;
        RECT 18.990 120.890 19.190 121.740 ;
        RECT 20.990 120.890 21.190 121.740 ;
        RECT 22.990 120.890 23.190 121.740 ;
        RECT 24.990 120.890 25.190 121.740 ;
        RECT 26.990 120.890 27.190 121.740 ;
        RECT 28.990 120.890 29.190 121.740 ;
        RECT 30.990 120.890 31.190 121.740 ;
        RECT 32.990 120.890 33.190 121.740 ;
        RECT 34.990 120.890 35.190 121.740 ;
        RECT 36.990 120.890 37.190 121.740 ;
        RECT 38.990 120.890 39.190 121.740 ;
        RECT 40.990 120.890 41.190 121.740 ;
        RECT 42.990 120.890 43.190 121.740 ;
        RECT 44.990 120.890 45.190 121.740 ;
        RECT 46.990 120.890 47.190 121.740 ;
        RECT 48.990 120.890 49.190 121.740 ;
        RECT 50.990 120.890 51.190 121.740 ;
        RECT 52.990 120.890 53.190 121.740 ;
        RECT 54.990 120.890 55.190 121.740 ;
        RECT 56.990 120.890 57.190 121.740 ;
        RECT 58.990 120.890 59.190 121.740 ;
        RECT 60.990 120.890 61.190 121.740 ;
        RECT 62.990 120.890 63.190 121.740 ;
        RECT 64.990 120.890 65.190 121.740 ;
        RECT 66.990 120.890 67.190 121.740 ;
        RECT 68.990 120.890 69.190 121.740 ;
        RECT 70.990 120.890 71.190 121.740 ;
        RECT 89.925 120.890 90.125 121.740 ;
        RECT 91.925 120.890 92.125 121.740 ;
        RECT 93.925 120.890 94.125 121.740 ;
        RECT 95.925 120.890 96.125 121.740 ;
        RECT 97.925 120.890 98.125 121.740 ;
        RECT 99.925 120.890 100.125 121.740 ;
        RECT 101.925 120.890 102.125 121.740 ;
        RECT 103.925 120.890 104.125 121.740 ;
        RECT 105.925 120.890 106.125 121.740 ;
        RECT 107.925 120.890 108.125 121.740 ;
        RECT 109.925 120.890 110.125 121.740 ;
        RECT 111.925 120.890 112.125 121.740 ;
        RECT 113.925 120.890 114.125 121.740 ;
        RECT 115.925 120.890 116.125 121.740 ;
        RECT 117.925 120.890 118.125 121.740 ;
        RECT 119.925 120.890 120.125 121.740 ;
        RECT 121.925 120.890 122.125 121.740 ;
        RECT 123.925 120.890 124.125 121.740 ;
        RECT 125.925 120.890 126.125 121.740 ;
        RECT 127.925 120.890 128.125 121.740 ;
        RECT 129.925 120.890 130.125 121.740 ;
        RECT 131.925 120.890 132.125 121.740 ;
        RECT 133.925 120.890 134.125 121.740 ;
        RECT 135.925 120.890 136.125 121.740 ;
        RECT 137.925 120.890 138.125 121.740 ;
        RECT 139.925 120.890 140.125 121.740 ;
        RECT 141.925 120.890 142.125 121.740 ;
        RECT 143.925 120.890 144.125 121.740 ;
        RECT 145.925 120.890 146.125 121.740 ;
        RECT 147.925 120.890 148.125 121.740 ;
        RECT 149.925 120.890 150.125 121.740 ;
        RECT 151.925 120.890 152.125 121.740 ;
        RECT 153.895 120.890 154.155 121.740 ;
        RECT 6.890 120.490 7.290 120.890 ;
        RECT 8.890 120.490 9.290 120.890 ;
        RECT 10.890 120.490 11.290 120.890 ;
        RECT 12.890 120.490 13.290 120.890 ;
        RECT 14.890 120.490 15.290 120.890 ;
        RECT 16.890 120.490 17.290 120.890 ;
        RECT 18.890 120.490 19.290 120.890 ;
        RECT 20.890 120.490 21.290 120.890 ;
        RECT 22.890 120.490 23.290 120.890 ;
        RECT 24.890 120.490 25.290 120.890 ;
        RECT 26.890 120.490 27.290 120.890 ;
        RECT 28.890 120.490 29.290 120.890 ;
        RECT 30.890 120.490 31.290 120.890 ;
        RECT 32.890 120.490 33.290 120.890 ;
        RECT 34.890 120.490 35.290 120.890 ;
        RECT 36.890 120.490 37.290 120.890 ;
        RECT 38.890 120.490 39.290 120.890 ;
        RECT 40.890 120.490 41.290 120.890 ;
        RECT 42.890 120.490 43.290 120.890 ;
        RECT 44.890 120.490 45.290 120.890 ;
        RECT 46.890 120.490 47.290 120.890 ;
        RECT 48.890 120.490 49.290 120.890 ;
        RECT 50.890 120.490 51.290 120.890 ;
        RECT 52.890 120.490 53.290 120.890 ;
        RECT 54.890 120.490 55.290 120.890 ;
        RECT 56.890 120.490 57.290 120.890 ;
        RECT 58.890 120.490 59.290 120.890 ;
        RECT 60.890 120.490 61.290 120.890 ;
        RECT 62.890 120.490 63.290 120.890 ;
        RECT 64.890 120.490 65.290 120.890 ;
        RECT 66.890 120.490 67.290 120.890 ;
        RECT 68.890 120.490 69.290 120.890 ;
        RECT 70.890 120.490 71.290 120.890 ;
        RECT 72.890 120.490 73.290 120.890 ;
        RECT 87.825 120.490 88.225 120.890 ;
        RECT 89.825 120.490 90.225 120.890 ;
        RECT 91.825 120.490 92.225 120.890 ;
        RECT 93.825 120.490 94.225 120.890 ;
        RECT 95.825 120.490 96.225 120.890 ;
        RECT 97.825 120.490 98.225 120.890 ;
        RECT 99.825 120.490 100.225 120.890 ;
        RECT 101.825 120.490 102.225 120.890 ;
        RECT 103.825 120.490 104.225 120.890 ;
        RECT 105.825 120.490 106.225 120.890 ;
        RECT 107.825 120.490 108.225 120.890 ;
        RECT 109.825 120.490 110.225 120.890 ;
        RECT 111.825 120.490 112.225 120.890 ;
        RECT 113.825 120.490 114.225 120.890 ;
        RECT 115.825 120.490 116.225 120.890 ;
        RECT 117.825 120.490 118.225 120.890 ;
        RECT 119.825 120.490 120.225 120.890 ;
        RECT 121.825 120.490 122.225 120.890 ;
        RECT 123.825 120.490 124.225 120.890 ;
        RECT 125.825 120.490 126.225 120.890 ;
        RECT 127.825 120.490 128.225 120.890 ;
        RECT 129.825 120.490 130.225 120.890 ;
        RECT 131.825 120.490 132.225 120.890 ;
        RECT 133.825 120.490 134.225 120.890 ;
        RECT 135.825 120.490 136.225 120.890 ;
        RECT 137.825 120.490 138.225 120.890 ;
        RECT 139.825 120.490 140.225 120.890 ;
        RECT 141.825 120.490 142.225 120.890 ;
        RECT 143.825 120.490 144.225 120.890 ;
        RECT 145.825 120.490 146.225 120.890 ;
        RECT 147.825 120.490 148.225 120.890 ;
        RECT 149.825 120.490 150.225 120.890 ;
        RECT 151.825 120.490 152.225 120.890 ;
        RECT 153.825 120.490 154.225 120.890 ;
        RECT 6.890 120.290 8.540 120.490 ;
        RECT 8.890 120.290 74.540 120.490 ;
        RECT 86.575 120.290 152.225 120.490 ;
        RECT 152.575 120.290 154.225 120.490 ;
        RECT 6.890 119.890 7.290 120.290 ;
        RECT 8.890 119.890 9.290 120.290 ;
        RECT 10.890 119.890 11.290 120.290 ;
        RECT 12.890 119.890 13.290 120.290 ;
        RECT 14.890 119.890 15.290 120.290 ;
        RECT 16.890 119.890 17.290 120.290 ;
        RECT 18.890 119.890 19.290 120.290 ;
        RECT 20.890 119.890 21.290 120.290 ;
        RECT 22.890 119.890 23.290 120.290 ;
        RECT 24.890 119.890 25.290 120.290 ;
        RECT 26.890 119.890 27.290 120.290 ;
        RECT 28.890 119.890 29.290 120.290 ;
        RECT 30.890 119.890 31.290 120.290 ;
        RECT 32.890 119.890 33.290 120.290 ;
        RECT 34.890 119.890 35.290 120.290 ;
        RECT 36.890 119.890 37.290 120.290 ;
        RECT 38.890 119.890 39.290 120.290 ;
        RECT 40.890 119.890 41.290 120.290 ;
        RECT 42.890 119.890 43.290 120.290 ;
        RECT 44.890 119.890 45.290 120.290 ;
        RECT 46.890 119.890 47.290 120.290 ;
        RECT 48.890 119.890 49.290 120.290 ;
        RECT 50.890 119.890 51.290 120.290 ;
        RECT 52.890 119.890 53.290 120.290 ;
        RECT 54.890 119.890 55.290 120.290 ;
        RECT 56.890 119.890 57.290 120.290 ;
        RECT 58.890 119.890 59.290 120.290 ;
        RECT 60.890 119.890 61.290 120.290 ;
        RECT 62.890 119.890 63.290 120.290 ;
        RECT 64.890 119.890 65.290 120.290 ;
        RECT 66.890 119.890 67.290 120.290 ;
        RECT 68.890 119.890 69.290 120.290 ;
        RECT 70.890 119.890 71.290 120.290 ;
        RECT 72.890 119.890 73.290 120.290 ;
        RECT 87.825 119.890 88.225 120.290 ;
        RECT 89.825 119.890 90.225 120.290 ;
        RECT 91.825 119.890 92.225 120.290 ;
        RECT 93.825 119.890 94.225 120.290 ;
        RECT 95.825 119.890 96.225 120.290 ;
        RECT 97.825 119.890 98.225 120.290 ;
        RECT 99.825 119.890 100.225 120.290 ;
        RECT 101.825 119.890 102.225 120.290 ;
        RECT 103.825 119.890 104.225 120.290 ;
        RECT 105.825 119.890 106.225 120.290 ;
        RECT 107.825 119.890 108.225 120.290 ;
        RECT 109.825 119.890 110.225 120.290 ;
        RECT 111.825 119.890 112.225 120.290 ;
        RECT 113.825 119.890 114.225 120.290 ;
        RECT 115.825 119.890 116.225 120.290 ;
        RECT 117.825 119.890 118.225 120.290 ;
        RECT 119.825 119.890 120.225 120.290 ;
        RECT 121.825 119.890 122.225 120.290 ;
        RECT 123.825 119.890 124.225 120.290 ;
        RECT 125.825 119.890 126.225 120.290 ;
        RECT 127.825 119.890 128.225 120.290 ;
        RECT 129.825 119.890 130.225 120.290 ;
        RECT 131.825 119.890 132.225 120.290 ;
        RECT 133.825 119.890 134.225 120.290 ;
        RECT 135.825 119.890 136.225 120.290 ;
        RECT 137.825 119.890 138.225 120.290 ;
        RECT 139.825 119.890 140.225 120.290 ;
        RECT 141.825 119.890 142.225 120.290 ;
        RECT 143.825 119.890 144.225 120.290 ;
        RECT 145.825 119.890 146.225 120.290 ;
        RECT 147.825 119.890 148.225 120.290 ;
        RECT 149.825 119.890 150.225 120.290 ;
        RECT 151.825 119.890 152.225 120.290 ;
        RECT 153.825 119.890 154.225 120.290 ;
        RECT 6.960 119.040 7.220 119.890 ;
        RECT 8.990 119.040 9.190 119.890 ;
        RECT 10.990 119.040 11.190 119.890 ;
        RECT 12.990 119.040 13.190 119.890 ;
        RECT 14.990 119.040 15.190 119.890 ;
        RECT 16.990 119.040 17.190 119.890 ;
        RECT 18.990 119.040 19.190 119.890 ;
        RECT 20.990 119.040 21.190 119.890 ;
        RECT 22.990 119.040 23.190 119.890 ;
        RECT 24.990 119.040 25.190 119.890 ;
        RECT 26.990 119.040 27.190 119.890 ;
        RECT 28.990 119.040 29.190 119.890 ;
        RECT 30.990 119.040 31.190 119.890 ;
        RECT 32.990 119.040 33.190 119.890 ;
        RECT 34.990 119.040 35.190 119.890 ;
        RECT 36.990 119.040 37.190 119.890 ;
        RECT 38.990 119.040 39.190 119.890 ;
        RECT 40.990 119.040 41.190 119.890 ;
        RECT 42.990 119.040 43.190 119.890 ;
        RECT 44.990 119.040 45.190 119.890 ;
        RECT 46.990 119.040 47.190 119.890 ;
        RECT 48.990 119.040 49.190 119.890 ;
        RECT 50.990 119.040 51.190 119.890 ;
        RECT 52.990 119.040 53.190 119.890 ;
        RECT 54.990 119.040 55.190 119.890 ;
        RECT 56.990 119.040 57.190 119.890 ;
        RECT 58.990 119.040 59.190 119.890 ;
        RECT 60.990 119.040 61.190 119.890 ;
        RECT 62.990 119.040 63.190 119.890 ;
        RECT 64.990 119.040 65.190 119.890 ;
        RECT 66.990 119.040 67.190 119.890 ;
        RECT 68.990 119.040 69.190 119.890 ;
        RECT 70.990 119.040 71.190 119.890 ;
        RECT 89.925 119.040 90.125 119.890 ;
        RECT 91.925 119.040 92.125 119.890 ;
        RECT 93.925 119.040 94.125 119.890 ;
        RECT 95.925 119.040 96.125 119.890 ;
        RECT 97.925 119.040 98.125 119.890 ;
        RECT 99.925 119.040 100.125 119.890 ;
        RECT 101.925 119.040 102.125 119.890 ;
        RECT 103.925 119.040 104.125 119.890 ;
        RECT 105.925 119.040 106.125 119.890 ;
        RECT 107.925 119.040 108.125 119.890 ;
        RECT 109.925 119.040 110.125 119.890 ;
        RECT 111.925 119.040 112.125 119.890 ;
        RECT 113.925 119.040 114.125 119.890 ;
        RECT 115.925 119.040 116.125 119.890 ;
        RECT 117.925 119.040 118.125 119.890 ;
        RECT 119.925 119.040 120.125 119.890 ;
        RECT 121.925 119.040 122.125 119.890 ;
        RECT 123.925 119.040 124.125 119.890 ;
        RECT 125.925 119.040 126.125 119.890 ;
        RECT 127.925 119.040 128.125 119.890 ;
        RECT 129.925 119.040 130.125 119.890 ;
        RECT 131.925 119.040 132.125 119.890 ;
        RECT 133.925 119.040 134.125 119.890 ;
        RECT 135.925 119.040 136.125 119.890 ;
        RECT 137.925 119.040 138.125 119.890 ;
        RECT 139.925 119.040 140.125 119.890 ;
        RECT 141.925 119.040 142.125 119.890 ;
        RECT 143.925 119.040 144.125 119.890 ;
        RECT 145.925 119.040 146.125 119.890 ;
        RECT 147.925 119.040 148.125 119.890 ;
        RECT 149.925 119.040 150.125 119.890 ;
        RECT 151.925 119.040 152.125 119.890 ;
        RECT 153.895 119.040 154.155 119.890 ;
        RECT 6.890 118.640 7.290 119.040 ;
        RECT 8.890 118.640 9.290 119.040 ;
        RECT 10.890 118.640 11.290 119.040 ;
        RECT 12.890 118.640 13.290 119.040 ;
        RECT 14.890 118.640 15.290 119.040 ;
        RECT 16.890 118.640 17.290 119.040 ;
        RECT 18.890 118.640 19.290 119.040 ;
        RECT 20.890 118.640 21.290 119.040 ;
        RECT 22.890 118.640 23.290 119.040 ;
        RECT 24.890 118.640 25.290 119.040 ;
        RECT 26.890 118.640 27.290 119.040 ;
        RECT 28.890 118.640 29.290 119.040 ;
        RECT 30.890 118.640 31.290 119.040 ;
        RECT 32.890 118.640 33.290 119.040 ;
        RECT 34.890 118.640 35.290 119.040 ;
        RECT 36.890 118.640 37.290 119.040 ;
        RECT 38.890 118.640 39.290 119.040 ;
        RECT 40.890 118.640 41.290 119.040 ;
        RECT 42.890 118.640 43.290 119.040 ;
        RECT 44.890 118.640 45.290 119.040 ;
        RECT 46.890 118.640 47.290 119.040 ;
        RECT 48.890 118.640 49.290 119.040 ;
        RECT 50.890 118.640 51.290 119.040 ;
        RECT 52.890 118.640 53.290 119.040 ;
        RECT 54.890 118.640 55.290 119.040 ;
        RECT 56.890 118.640 57.290 119.040 ;
        RECT 58.890 118.640 59.290 119.040 ;
        RECT 60.890 118.640 61.290 119.040 ;
        RECT 62.890 118.640 63.290 119.040 ;
        RECT 64.890 118.640 65.290 119.040 ;
        RECT 66.890 118.640 67.290 119.040 ;
        RECT 68.890 118.640 69.290 119.040 ;
        RECT 70.890 118.640 71.290 119.040 ;
        RECT 72.890 118.640 73.290 119.040 ;
        RECT 87.825 118.640 88.225 119.040 ;
        RECT 89.825 118.640 90.225 119.040 ;
        RECT 91.825 118.640 92.225 119.040 ;
        RECT 93.825 118.640 94.225 119.040 ;
        RECT 95.825 118.640 96.225 119.040 ;
        RECT 97.825 118.640 98.225 119.040 ;
        RECT 99.825 118.640 100.225 119.040 ;
        RECT 101.825 118.640 102.225 119.040 ;
        RECT 103.825 118.640 104.225 119.040 ;
        RECT 105.825 118.640 106.225 119.040 ;
        RECT 107.825 118.640 108.225 119.040 ;
        RECT 109.825 118.640 110.225 119.040 ;
        RECT 111.825 118.640 112.225 119.040 ;
        RECT 113.825 118.640 114.225 119.040 ;
        RECT 115.825 118.640 116.225 119.040 ;
        RECT 117.825 118.640 118.225 119.040 ;
        RECT 119.825 118.640 120.225 119.040 ;
        RECT 121.825 118.640 122.225 119.040 ;
        RECT 123.825 118.640 124.225 119.040 ;
        RECT 125.825 118.640 126.225 119.040 ;
        RECT 127.825 118.640 128.225 119.040 ;
        RECT 129.825 118.640 130.225 119.040 ;
        RECT 131.825 118.640 132.225 119.040 ;
        RECT 133.825 118.640 134.225 119.040 ;
        RECT 135.825 118.640 136.225 119.040 ;
        RECT 137.825 118.640 138.225 119.040 ;
        RECT 139.825 118.640 140.225 119.040 ;
        RECT 141.825 118.640 142.225 119.040 ;
        RECT 143.825 118.640 144.225 119.040 ;
        RECT 145.825 118.640 146.225 119.040 ;
        RECT 147.825 118.640 148.225 119.040 ;
        RECT 149.825 118.640 150.225 119.040 ;
        RECT 151.825 118.640 152.225 119.040 ;
        RECT 153.825 118.640 154.225 119.040 ;
        RECT 6.890 118.440 8.540 118.640 ;
        RECT 8.890 118.440 74.540 118.640 ;
        RECT 86.575 118.440 152.225 118.640 ;
        RECT 152.575 118.440 154.225 118.640 ;
        RECT 6.890 118.040 7.290 118.440 ;
        RECT 8.890 118.040 9.290 118.440 ;
        RECT 10.890 118.040 11.290 118.440 ;
        RECT 12.890 118.040 13.290 118.440 ;
        RECT 14.890 118.040 15.290 118.440 ;
        RECT 16.890 118.040 17.290 118.440 ;
        RECT 18.890 118.040 19.290 118.440 ;
        RECT 20.890 118.040 21.290 118.440 ;
        RECT 22.890 118.040 23.290 118.440 ;
        RECT 24.890 118.040 25.290 118.440 ;
        RECT 26.890 118.040 27.290 118.440 ;
        RECT 28.890 118.040 29.290 118.440 ;
        RECT 30.890 118.040 31.290 118.440 ;
        RECT 32.890 118.040 33.290 118.440 ;
        RECT 34.890 118.040 35.290 118.440 ;
        RECT 36.890 118.040 37.290 118.440 ;
        RECT 38.890 118.040 39.290 118.440 ;
        RECT 40.890 118.040 41.290 118.440 ;
        RECT 42.890 118.040 43.290 118.440 ;
        RECT 44.890 118.040 45.290 118.440 ;
        RECT 46.890 118.040 47.290 118.440 ;
        RECT 48.890 118.040 49.290 118.440 ;
        RECT 50.890 118.040 51.290 118.440 ;
        RECT 52.890 118.040 53.290 118.440 ;
        RECT 54.890 118.040 55.290 118.440 ;
        RECT 56.890 118.040 57.290 118.440 ;
        RECT 58.890 118.040 59.290 118.440 ;
        RECT 60.890 118.040 61.290 118.440 ;
        RECT 62.890 118.040 63.290 118.440 ;
        RECT 64.890 118.040 65.290 118.440 ;
        RECT 66.890 118.040 67.290 118.440 ;
        RECT 68.890 118.040 69.290 118.440 ;
        RECT 70.890 118.040 71.290 118.440 ;
        RECT 72.890 118.040 73.290 118.440 ;
        RECT 87.825 118.040 88.225 118.440 ;
        RECT 89.825 118.040 90.225 118.440 ;
        RECT 91.825 118.040 92.225 118.440 ;
        RECT 93.825 118.040 94.225 118.440 ;
        RECT 95.825 118.040 96.225 118.440 ;
        RECT 97.825 118.040 98.225 118.440 ;
        RECT 99.825 118.040 100.225 118.440 ;
        RECT 101.825 118.040 102.225 118.440 ;
        RECT 103.825 118.040 104.225 118.440 ;
        RECT 105.825 118.040 106.225 118.440 ;
        RECT 107.825 118.040 108.225 118.440 ;
        RECT 109.825 118.040 110.225 118.440 ;
        RECT 111.825 118.040 112.225 118.440 ;
        RECT 113.825 118.040 114.225 118.440 ;
        RECT 115.825 118.040 116.225 118.440 ;
        RECT 117.825 118.040 118.225 118.440 ;
        RECT 119.825 118.040 120.225 118.440 ;
        RECT 121.825 118.040 122.225 118.440 ;
        RECT 123.825 118.040 124.225 118.440 ;
        RECT 125.825 118.040 126.225 118.440 ;
        RECT 127.825 118.040 128.225 118.440 ;
        RECT 129.825 118.040 130.225 118.440 ;
        RECT 131.825 118.040 132.225 118.440 ;
        RECT 133.825 118.040 134.225 118.440 ;
        RECT 135.825 118.040 136.225 118.440 ;
        RECT 137.825 118.040 138.225 118.440 ;
        RECT 139.825 118.040 140.225 118.440 ;
        RECT 141.825 118.040 142.225 118.440 ;
        RECT 143.825 118.040 144.225 118.440 ;
        RECT 145.825 118.040 146.225 118.440 ;
        RECT 147.825 118.040 148.225 118.440 ;
        RECT 149.825 118.040 150.225 118.440 ;
        RECT 151.825 118.040 152.225 118.440 ;
        RECT 153.825 118.040 154.225 118.440 ;
        RECT 6.960 117.190 7.220 118.040 ;
        RECT 8.990 117.190 9.190 118.040 ;
        RECT 10.990 117.190 11.190 118.040 ;
        RECT 12.990 117.190 13.190 118.040 ;
        RECT 14.990 117.190 15.190 118.040 ;
        RECT 16.990 117.190 17.190 118.040 ;
        RECT 18.990 117.190 19.190 118.040 ;
        RECT 20.990 117.190 21.190 118.040 ;
        RECT 22.990 117.190 23.190 118.040 ;
        RECT 24.990 117.190 25.190 118.040 ;
        RECT 26.990 117.190 27.190 118.040 ;
        RECT 28.990 117.190 29.190 118.040 ;
        RECT 30.990 117.190 31.190 118.040 ;
        RECT 32.990 117.190 33.190 118.040 ;
        RECT 34.990 117.190 35.190 118.040 ;
        RECT 36.990 117.190 37.190 118.040 ;
        RECT 38.990 117.190 39.190 118.040 ;
        RECT 40.990 117.190 41.190 118.040 ;
        RECT 42.990 117.190 43.190 118.040 ;
        RECT 44.990 117.190 45.190 118.040 ;
        RECT 46.990 117.190 47.190 118.040 ;
        RECT 48.990 117.190 49.190 118.040 ;
        RECT 50.990 117.190 51.190 118.040 ;
        RECT 52.990 117.190 53.190 118.040 ;
        RECT 54.990 117.190 55.190 118.040 ;
        RECT 56.990 117.190 57.190 118.040 ;
        RECT 58.990 117.190 59.190 118.040 ;
        RECT 60.990 117.190 61.190 118.040 ;
        RECT 62.990 117.190 63.190 118.040 ;
        RECT 64.990 117.190 65.190 118.040 ;
        RECT 66.990 117.190 67.190 118.040 ;
        RECT 68.990 117.190 69.190 118.040 ;
        RECT 70.990 117.190 71.190 118.040 ;
        RECT 89.925 117.190 90.125 118.040 ;
        RECT 91.925 117.190 92.125 118.040 ;
        RECT 93.925 117.190 94.125 118.040 ;
        RECT 95.925 117.190 96.125 118.040 ;
        RECT 97.925 117.190 98.125 118.040 ;
        RECT 99.925 117.190 100.125 118.040 ;
        RECT 101.925 117.190 102.125 118.040 ;
        RECT 103.925 117.190 104.125 118.040 ;
        RECT 105.925 117.190 106.125 118.040 ;
        RECT 107.925 117.190 108.125 118.040 ;
        RECT 109.925 117.190 110.125 118.040 ;
        RECT 111.925 117.190 112.125 118.040 ;
        RECT 113.925 117.190 114.125 118.040 ;
        RECT 115.925 117.190 116.125 118.040 ;
        RECT 117.925 117.190 118.125 118.040 ;
        RECT 119.925 117.190 120.125 118.040 ;
        RECT 121.925 117.190 122.125 118.040 ;
        RECT 123.925 117.190 124.125 118.040 ;
        RECT 125.925 117.190 126.125 118.040 ;
        RECT 127.925 117.190 128.125 118.040 ;
        RECT 129.925 117.190 130.125 118.040 ;
        RECT 131.925 117.190 132.125 118.040 ;
        RECT 133.925 117.190 134.125 118.040 ;
        RECT 135.925 117.190 136.125 118.040 ;
        RECT 137.925 117.190 138.125 118.040 ;
        RECT 139.925 117.190 140.125 118.040 ;
        RECT 141.925 117.190 142.125 118.040 ;
        RECT 143.925 117.190 144.125 118.040 ;
        RECT 145.925 117.190 146.125 118.040 ;
        RECT 147.925 117.190 148.125 118.040 ;
        RECT 149.925 117.190 150.125 118.040 ;
        RECT 151.925 117.190 152.125 118.040 ;
        RECT 153.895 117.190 154.155 118.040 ;
        RECT 6.890 116.790 7.290 117.190 ;
        RECT 8.890 116.790 9.290 117.190 ;
        RECT 10.890 116.790 11.290 117.190 ;
        RECT 12.890 116.790 13.290 117.190 ;
        RECT 14.890 116.790 15.290 117.190 ;
        RECT 16.890 116.790 17.290 117.190 ;
        RECT 18.890 116.790 19.290 117.190 ;
        RECT 20.890 116.790 21.290 117.190 ;
        RECT 22.890 116.790 23.290 117.190 ;
        RECT 24.890 116.790 25.290 117.190 ;
        RECT 26.890 116.790 27.290 117.190 ;
        RECT 28.890 116.790 29.290 117.190 ;
        RECT 30.890 116.790 31.290 117.190 ;
        RECT 32.890 116.790 33.290 117.190 ;
        RECT 34.890 116.790 35.290 117.190 ;
        RECT 36.890 116.790 37.290 117.190 ;
        RECT 38.890 116.790 39.290 117.190 ;
        RECT 40.890 116.790 41.290 117.190 ;
        RECT 42.890 116.790 43.290 117.190 ;
        RECT 44.890 116.790 45.290 117.190 ;
        RECT 46.890 116.790 47.290 117.190 ;
        RECT 48.890 116.790 49.290 117.190 ;
        RECT 50.890 116.790 51.290 117.190 ;
        RECT 52.890 116.790 53.290 117.190 ;
        RECT 54.890 116.790 55.290 117.190 ;
        RECT 56.890 116.790 57.290 117.190 ;
        RECT 58.890 116.790 59.290 117.190 ;
        RECT 60.890 116.790 61.290 117.190 ;
        RECT 62.890 116.790 63.290 117.190 ;
        RECT 64.890 116.790 65.290 117.190 ;
        RECT 66.890 116.790 67.290 117.190 ;
        RECT 68.890 116.790 69.290 117.190 ;
        RECT 70.890 116.790 71.290 117.190 ;
        RECT 72.890 116.790 73.290 117.190 ;
        RECT 87.825 116.790 88.225 117.190 ;
        RECT 89.825 116.790 90.225 117.190 ;
        RECT 91.825 116.790 92.225 117.190 ;
        RECT 93.825 116.790 94.225 117.190 ;
        RECT 95.825 116.790 96.225 117.190 ;
        RECT 97.825 116.790 98.225 117.190 ;
        RECT 99.825 116.790 100.225 117.190 ;
        RECT 101.825 116.790 102.225 117.190 ;
        RECT 103.825 116.790 104.225 117.190 ;
        RECT 105.825 116.790 106.225 117.190 ;
        RECT 107.825 116.790 108.225 117.190 ;
        RECT 109.825 116.790 110.225 117.190 ;
        RECT 111.825 116.790 112.225 117.190 ;
        RECT 113.825 116.790 114.225 117.190 ;
        RECT 115.825 116.790 116.225 117.190 ;
        RECT 117.825 116.790 118.225 117.190 ;
        RECT 119.825 116.790 120.225 117.190 ;
        RECT 121.825 116.790 122.225 117.190 ;
        RECT 123.825 116.790 124.225 117.190 ;
        RECT 125.825 116.790 126.225 117.190 ;
        RECT 127.825 116.790 128.225 117.190 ;
        RECT 129.825 116.790 130.225 117.190 ;
        RECT 131.825 116.790 132.225 117.190 ;
        RECT 133.825 116.790 134.225 117.190 ;
        RECT 135.825 116.790 136.225 117.190 ;
        RECT 137.825 116.790 138.225 117.190 ;
        RECT 139.825 116.790 140.225 117.190 ;
        RECT 141.825 116.790 142.225 117.190 ;
        RECT 143.825 116.790 144.225 117.190 ;
        RECT 145.825 116.790 146.225 117.190 ;
        RECT 147.825 116.790 148.225 117.190 ;
        RECT 149.825 116.790 150.225 117.190 ;
        RECT 151.825 116.790 152.225 117.190 ;
        RECT 153.825 116.790 154.225 117.190 ;
        RECT 6.890 116.590 8.540 116.790 ;
        RECT 8.890 116.590 74.540 116.790 ;
        RECT 86.575 116.590 152.225 116.790 ;
        RECT 152.575 116.590 154.225 116.790 ;
        RECT 6.890 116.190 7.290 116.590 ;
        RECT 8.890 116.190 9.290 116.590 ;
        RECT 10.890 116.190 11.290 116.590 ;
        RECT 12.890 116.190 13.290 116.590 ;
        RECT 14.890 116.190 15.290 116.590 ;
        RECT 16.890 116.190 17.290 116.590 ;
        RECT 18.890 116.190 19.290 116.590 ;
        RECT 20.890 116.190 21.290 116.590 ;
        RECT 22.890 116.190 23.290 116.590 ;
        RECT 24.890 116.190 25.290 116.590 ;
        RECT 26.890 116.190 27.290 116.590 ;
        RECT 28.890 116.190 29.290 116.590 ;
        RECT 30.890 116.190 31.290 116.590 ;
        RECT 32.890 116.190 33.290 116.590 ;
        RECT 34.890 116.190 35.290 116.590 ;
        RECT 36.890 116.190 37.290 116.590 ;
        RECT 38.890 116.190 39.290 116.590 ;
        RECT 40.890 116.190 41.290 116.590 ;
        RECT 42.890 116.190 43.290 116.590 ;
        RECT 44.890 116.190 45.290 116.590 ;
        RECT 46.890 116.190 47.290 116.590 ;
        RECT 48.890 116.190 49.290 116.590 ;
        RECT 50.890 116.190 51.290 116.590 ;
        RECT 52.890 116.190 53.290 116.590 ;
        RECT 54.890 116.190 55.290 116.590 ;
        RECT 56.890 116.190 57.290 116.590 ;
        RECT 58.890 116.190 59.290 116.590 ;
        RECT 60.890 116.190 61.290 116.590 ;
        RECT 62.890 116.190 63.290 116.590 ;
        RECT 64.890 116.190 65.290 116.590 ;
        RECT 66.890 116.190 67.290 116.590 ;
        RECT 68.890 116.190 69.290 116.590 ;
        RECT 70.890 116.190 71.290 116.590 ;
        RECT 72.890 116.190 73.290 116.590 ;
        RECT 87.825 116.190 88.225 116.590 ;
        RECT 89.825 116.190 90.225 116.590 ;
        RECT 91.825 116.190 92.225 116.590 ;
        RECT 93.825 116.190 94.225 116.590 ;
        RECT 95.825 116.190 96.225 116.590 ;
        RECT 97.825 116.190 98.225 116.590 ;
        RECT 99.825 116.190 100.225 116.590 ;
        RECT 101.825 116.190 102.225 116.590 ;
        RECT 103.825 116.190 104.225 116.590 ;
        RECT 105.825 116.190 106.225 116.590 ;
        RECT 107.825 116.190 108.225 116.590 ;
        RECT 109.825 116.190 110.225 116.590 ;
        RECT 111.825 116.190 112.225 116.590 ;
        RECT 113.825 116.190 114.225 116.590 ;
        RECT 115.825 116.190 116.225 116.590 ;
        RECT 117.825 116.190 118.225 116.590 ;
        RECT 119.825 116.190 120.225 116.590 ;
        RECT 121.825 116.190 122.225 116.590 ;
        RECT 123.825 116.190 124.225 116.590 ;
        RECT 125.825 116.190 126.225 116.590 ;
        RECT 127.825 116.190 128.225 116.590 ;
        RECT 129.825 116.190 130.225 116.590 ;
        RECT 131.825 116.190 132.225 116.590 ;
        RECT 133.825 116.190 134.225 116.590 ;
        RECT 135.825 116.190 136.225 116.590 ;
        RECT 137.825 116.190 138.225 116.590 ;
        RECT 139.825 116.190 140.225 116.590 ;
        RECT 141.825 116.190 142.225 116.590 ;
        RECT 143.825 116.190 144.225 116.590 ;
        RECT 145.825 116.190 146.225 116.590 ;
        RECT 147.825 116.190 148.225 116.590 ;
        RECT 149.825 116.190 150.225 116.590 ;
        RECT 151.825 116.190 152.225 116.590 ;
        RECT 153.825 116.190 154.225 116.590 ;
        RECT 6.960 115.340 7.220 116.190 ;
        RECT 8.990 115.340 9.190 116.190 ;
        RECT 10.990 115.340 11.190 116.190 ;
        RECT 12.990 115.340 13.190 116.190 ;
        RECT 14.990 115.340 15.190 116.190 ;
        RECT 16.990 115.340 17.190 116.190 ;
        RECT 18.990 115.340 19.190 116.190 ;
        RECT 20.990 115.340 21.190 116.190 ;
        RECT 22.990 115.340 23.190 116.190 ;
        RECT 24.990 115.340 25.190 116.190 ;
        RECT 26.990 115.340 27.190 116.190 ;
        RECT 28.990 115.340 29.190 116.190 ;
        RECT 30.990 115.340 31.190 116.190 ;
        RECT 32.990 115.340 33.190 116.190 ;
        RECT 34.990 115.340 35.190 116.190 ;
        RECT 36.990 115.340 37.190 116.190 ;
        RECT 38.990 115.340 39.190 116.190 ;
        RECT 40.990 115.340 41.190 116.190 ;
        RECT 42.990 115.340 43.190 116.190 ;
        RECT 44.990 115.340 45.190 116.190 ;
        RECT 46.990 115.340 47.190 116.190 ;
        RECT 48.990 115.340 49.190 116.190 ;
        RECT 50.990 115.340 51.190 116.190 ;
        RECT 52.990 115.340 53.190 116.190 ;
        RECT 54.990 115.340 55.190 116.190 ;
        RECT 56.990 115.340 57.190 116.190 ;
        RECT 58.990 115.340 59.190 116.190 ;
        RECT 60.990 115.340 61.190 116.190 ;
        RECT 62.990 115.340 63.190 116.190 ;
        RECT 64.990 115.340 65.190 116.190 ;
        RECT 66.990 115.340 67.190 116.190 ;
        RECT 68.990 115.340 69.190 116.190 ;
        RECT 70.990 115.340 71.190 116.190 ;
        RECT 89.925 115.340 90.125 116.190 ;
        RECT 91.925 115.340 92.125 116.190 ;
        RECT 93.925 115.340 94.125 116.190 ;
        RECT 95.925 115.340 96.125 116.190 ;
        RECT 97.925 115.340 98.125 116.190 ;
        RECT 99.925 115.340 100.125 116.190 ;
        RECT 101.925 115.340 102.125 116.190 ;
        RECT 103.925 115.340 104.125 116.190 ;
        RECT 105.925 115.340 106.125 116.190 ;
        RECT 107.925 115.340 108.125 116.190 ;
        RECT 109.925 115.340 110.125 116.190 ;
        RECT 111.925 115.340 112.125 116.190 ;
        RECT 113.925 115.340 114.125 116.190 ;
        RECT 115.925 115.340 116.125 116.190 ;
        RECT 117.925 115.340 118.125 116.190 ;
        RECT 119.925 115.340 120.125 116.190 ;
        RECT 121.925 115.340 122.125 116.190 ;
        RECT 123.925 115.340 124.125 116.190 ;
        RECT 125.925 115.340 126.125 116.190 ;
        RECT 127.925 115.340 128.125 116.190 ;
        RECT 129.925 115.340 130.125 116.190 ;
        RECT 131.925 115.340 132.125 116.190 ;
        RECT 133.925 115.340 134.125 116.190 ;
        RECT 135.925 115.340 136.125 116.190 ;
        RECT 137.925 115.340 138.125 116.190 ;
        RECT 139.925 115.340 140.125 116.190 ;
        RECT 141.925 115.340 142.125 116.190 ;
        RECT 143.925 115.340 144.125 116.190 ;
        RECT 145.925 115.340 146.125 116.190 ;
        RECT 147.925 115.340 148.125 116.190 ;
        RECT 149.925 115.340 150.125 116.190 ;
        RECT 151.925 115.340 152.125 116.190 ;
        RECT 153.895 115.340 154.155 116.190 ;
        RECT 6.890 114.940 7.290 115.340 ;
        RECT 8.890 114.940 9.290 115.340 ;
        RECT 10.890 114.940 11.290 115.340 ;
        RECT 12.890 114.940 13.290 115.340 ;
        RECT 14.890 114.940 15.290 115.340 ;
        RECT 16.890 114.940 17.290 115.340 ;
        RECT 18.890 114.940 19.290 115.340 ;
        RECT 20.890 114.940 21.290 115.340 ;
        RECT 22.890 114.940 23.290 115.340 ;
        RECT 24.890 114.940 25.290 115.340 ;
        RECT 26.890 114.940 27.290 115.340 ;
        RECT 28.890 114.940 29.290 115.340 ;
        RECT 30.890 114.940 31.290 115.340 ;
        RECT 32.890 114.940 33.290 115.340 ;
        RECT 34.890 114.940 35.290 115.340 ;
        RECT 36.890 114.940 37.290 115.340 ;
        RECT 38.890 114.940 39.290 115.340 ;
        RECT 40.890 114.940 41.290 115.340 ;
        RECT 42.890 114.940 43.290 115.340 ;
        RECT 44.890 114.940 45.290 115.340 ;
        RECT 46.890 114.940 47.290 115.340 ;
        RECT 48.890 114.940 49.290 115.340 ;
        RECT 50.890 114.940 51.290 115.340 ;
        RECT 52.890 114.940 53.290 115.340 ;
        RECT 54.890 114.940 55.290 115.340 ;
        RECT 56.890 114.940 57.290 115.340 ;
        RECT 58.890 114.940 59.290 115.340 ;
        RECT 60.890 114.940 61.290 115.340 ;
        RECT 62.890 114.940 63.290 115.340 ;
        RECT 64.890 114.940 65.290 115.340 ;
        RECT 66.890 114.940 67.290 115.340 ;
        RECT 68.890 114.940 69.290 115.340 ;
        RECT 70.890 114.940 71.290 115.340 ;
        RECT 72.890 114.940 73.290 115.340 ;
        RECT 87.825 114.940 88.225 115.340 ;
        RECT 89.825 114.940 90.225 115.340 ;
        RECT 91.825 114.940 92.225 115.340 ;
        RECT 93.825 114.940 94.225 115.340 ;
        RECT 95.825 114.940 96.225 115.340 ;
        RECT 97.825 114.940 98.225 115.340 ;
        RECT 99.825 114.940 100.225 115.340 ;
        RECT 101.825 114.940 102.225 115.340 ;
        RECT 103.825 114.940 104.225 115.340 ;
        RECT 105.825 114.940 106.225 115.340 ;
        RECT 107.825 114.940 108.225 115.340 ;
        RECT 109.825 114.940 110.225 115.340 ;
        RECT 111.825 114.940 112.225 115.340 ;
        RECT 113.825 114.940 114.225 115.340 ;
        RECT 115.825 114.940 116.225 115.340 ;
        RECT 117.825 114.940 118.225 115.340 ;
        RECT 119.825 114.940 120.225 115.340 ;
        RECT 121.825 114.940 122.225 115.340 ;
        RECT 123.825 114.940 124.225 115.340 ;
        RECT 125.825 114.940 126.225 115.340 ;
        RECT 127.825 114.940 128.225 115.340 ;
        RECT 129.825 114.940 130.225 115.340 ;
        RECT 131.825 114.940 132.225 115.340 ;
        RECT 133.825 114.940 134.225 115.340 ;
        RECT 135.825 114.940 136.225 115.340 ;
        RECT 137.825 114.940 138.225 115.340 ;
        RECT 139.825 114.940 140.225 115.340 ;
        RECT 141.825 114.940 142.225 115.340 ;
        RECT 143.825 114.940 144.225 115.340 ;
        RECT 145.825 114.940 146.225 115.340 ;
        RECT 147.825 114.940 148.225 115.340 ;
        RECT 149.825 114.940 150.225 115.340 ;
        RECT 151.825 114.940 152.225 115.340 ;
        RECT 153.825 114.940 154.225 115.340 ;
        RECT 6.890 114.740 8.540 114.940 ;
        RECT 8.890 114.740 74.540 114.940 ;
        RECT 86.575 114.740 152.225 114.940 ;
        RECT 152.575 114.740 154.225 114.940 ;
        RECT 6.890 114.340 7.290 114.740 ;
        RECT 8.890 114.340 9.290 114.740 ;
        RECT 10.890 114.340 11.290 114.740 ;
        RECT 12.890 114.340 13.290 114.740 ;
        RECT 14.890 114.340 15.290 114.740 ;
        RECT 16.890 114.340 17.290 114.740 ;
        RECT 18.890 114.340 19.290 114.740 ;
        RECT 20.890 114.340 21.290 114.740 ;
        RECT 22.890 114.340 23.290 114.740 ;
        RECT 24.890 114.340 25.290 114.740 ;
        RECT 26.890 114.340 27.290 114.740 ;
        RECT 28.890 114.340 29.290 114.740 ;
        RECT 30.890 114.340 31.290 114.740 ;
        RECT 32.890 114.340 33.290 114.740 ;
        RECT 34.890 114.340 35.290 114.740 ;
        RECT 36.890 114.340 37.290 114.740 ;
        RECT 38.890 114.340 39.290 114.740 ;
        RECT 40.890 114.340 41.290 114.740 ;
        RECT 42.890 114.340 43.290 114.740 ;
        RECT 44.890 114.340 45.290 114.740 ;
        RECT 46.890 114.340 47.290 114.740 ;
        RECT 48.890 114.340 49.290 114.740 ;
        RECT 50.890 114.340 51.290 114.740 ;
        RECT 52.890 114.340 53.290 114.740 ;
        RECT 54.890 114.340 55.290 114.740 ;
        RECT 56.890 114.340 57.290 114.740 ;
        RECT 58.890 114.340 59.290 114.740 ;
        RECT 60.890 114.340 61.290 114.740 ;
        RECT 62.890 114.340 63.290 114.740 ;
        RECT 64.890 114.340 65.290 114.740 ;
        RECT 66.890 114.340 67.290 114.740 ;
        RECT 68.890 114.340 69.290 114.740 ;
        RECT 70.890 114.340 71.290 114.740 ;
        RECT 72.890 114.340 73.290 114.740 ;
        RECT 87.825 114.340 88.225 114.740 ;
        RECT 89.825 114.340 90.225 114.740 ;
        RECT 91.825 114.340 92.225 114.740 ;
        RECT 93.825 114.340 94.225 114.740 ;
        RECT 95.825 114.340 96.225 114.740 ;
        RECT 97.825 114.340 98.225 114.740 ;
        RECT 99.825 114.340 100.225 114.740 ;
        RECT 101.825 114.340 102.225 114.740 ;
        RECT 103.825 114.340 104.225 114.740 ;
        RECT 105.825 114.340 106.225 114.740 ;
        RECT 107.825 114.340 108.225 114.740 ;
        RECT 109.825 114.340 110.225 114.740 ;
        RECT 111.825 114.340 112.225 114.740 ;
        RECT 113.825 114.340 114.225 114.740 ;
        RECT 115.825 114.340 116.225 114.740 ;
        RECT 117.825 114.340 118.225 114.740 ;
        RECT 119.825 114.340 120.225 114.740 ;
        RECT 121.825 114.340 122.225 114.740 ;
        RECT 123.825 114.340 124.225 114.740 ;
        RECT 125.825 114.340 126.225 114.740 ;
        RECT 127.825 114.340 128.225 114.740 ;
        RECT 129.825 114.340 130.225 114.740 ;
        RECT 131.825 114.340 132.225 114.740 ;
        RECT 133.825 114.340 134.225 114.740 ;
        RECT 135.825 114.340 136.225 114.740 ;
        RECT 137.825 114.340 138.225 114.740 ;
        RECT 139.825 114.340 140.225 114.740 ;
        RECT 141.825 114.340 142.225 114.740 ;
        RECT 143.825 114.340 144.225 114.740 ;
        RECT 145.825 114.340 146.225 114.740 ;
        RECT 147.825 114.340 148.225 114.740 ;
        RECT 149.825 114.340 150.225 114.740 ;
        RECT 151.825 114.340 152.225 114.740 ;
        RECT 153.825 114.340 154.225 114.740 ;
        RECT 6.960 113.490 7.220 114.340 ;
        RECT 8.990 113.490 9.190 114.340 ;
        RECT 10.990 113.490 11.190 114.340 ;
        RECT 12.990 113.490 13.190 114.340 ;
        RECT 14.990 113.490 15.190 114.340 ;
        RECT 16.990 113.490 17.190 114.340 ;
        RECT 18.990 113.490 19.190 114.340 ;
        RECT 20.990 113.490 21.190 114.340 ;
        RECT 22.990 113.490 23.190 114.340 ;
        RECT 24.990 113.490 25.190 114.340 ;
        RECT 26.990 113.490 27.190 114.340 ;
        RECT 28.990 113.490 29.190 114.340 ;
        RECT 30.990 113.490 31.190 114.340 ;
        RECT 32.990 113.490 33.190 114.340 ;
        RECT 34.990 113.490 35.190 114.340 ;
        RECT 36.990 113.490 37.190 114.340 ;
        RECT 38.990 113.490 39.190 114.340 ;
        RECT 40.990 113.490 41.190 114.340 ;
        RECT 42.990 113.490 43.190 114.340 ;
        RECT 44.990 113.490 45.190 114.340 ;
        RECT 46.990 113.490 47.190 114.340 ;
        RECT 48.990 113.490 49.190 114.340 ;
        RECT 50.990 113.490 51.190 114.340 ;
        RECT 52.990 113.490 53.190 114.340 ;
        RECT 54.990 113.490 55.190 114.340 ;
        RECT 56.990 113.490 57.190 114.340 ;
        RECT 58.990 113.490 59.190 114.340 ;
        RECT 60.990 113.490 61.190 114.340 ;
        RECT 62.990 113.490 63.190 114.340 ;
        RECT 64.990 113.490 65.190 114.340 ;
        RECT 66.990 113.490 67.190 114.340 ;
        RECT 68.990 113.490 69.190 114.340 ;
        RECT 70.990 113.490 71.190 114.340 ;
        RECT 89.925 113.490 90.125 114.340 ;
        RECT 91.925 113.490 92.125 114.340 ;
        RECT 93.925 113.490 94.125 114.340 ;
        RECT 95.925 113.490 96.125 114.340 ;
        RECT 97.925 113.490 98.125 114.340 ;
        RECT 99.925 113.490 100.125 114.340 ;
        RECT 101.925 113.490 102.125 114.340 ;
        RECT 103.925 113.490 104.125 114.340 ;
        RECT 105.925 113.490 106.125 114.340 ;
        RECT 107.925 113.490 108.125 114.340 ;
        RECT 109.925 113.490 110.125 114.340 ;
        RECT 111.925 113.490 112.125 114.340 ;
        RECT 113.925 113.490 114.125 114.340 ;
        RECT 115.925 113.490 116.125 114.340 ;
        RECT 117.925 113.490 118.125 114.340 ;
        RECT 119.925 113.490 120.125 114.340 ;
        RECT 121.925 113.490 122.125 114.340 ;
        RECT 123.925 113.490 124.125 114.340 ;
        RECT 125.925 113.490 126.125 114.340 ;
        RECT 127.925 113.490 128.125 114.340 ;
        RECT 129.925 113.490 130.125 114.340 ;
        RECT 131.925 113.490 132.125 114.340 ;
        RECT 133.925 113.490 134.125 114.340 ;
        RECT 135.925 113.490 136.125 114.340 ;
        RECT 137.925 113.490 138.125 114.340 ;
        RECT 139.925 113.490 140.125 114.340 ;
        RECT 141.925 113.490 142.125 114.340 ;
        RECT 143.925 113.490 144.125 114.340 ;
        RECT 145.925 113.490 146.125 114.340 ;
        RECT 147.925 113.490 148.125 114.340 ;
        RECT 149.925 113.490 150.125 114.340 ;
        RECT 151.925 113.490 152.125 114.340 ;
        RECT 153.895 113.490 154.155 114.340 ;
        RECT 6.890 113.090 7.290 113.490 ;
        RECT 8.890 113.090 9.290 113.490 ;
        RECT 10.890 113.090 11.290 113.490 ;
        RECT 12.890 113.090 13.290 113.490 ;
        RECT 14.890 113.090 15.290 113.490 ;
        RECT 16.890 113.090 17.290 113.490 ;
        RECT 18.890 113.090 19.290 113.490 ;
        RECT 20.890 113.090 21.290 113.490 ;
        RECT 22.890 113.090 23.290 113.490 ;
        RECT 24.890 113.090 25.290 113.490 ;
        RECT 26.890 113.090 27.290 113.490 ;
        RECT 28.890 113.090 29.290 113.490 ;
        RECT 30.890 113.090 31.290 113.490 ;
        RECT 32.890 113.090 33.290 113.490 ;
        RECT 34.890 113.090 35.290 113.490 ;
        RECT 36.890 113.090 37.290 113.490 ;
        RECT 38.890 113.090 39.290 113.490 ;
        RECT 40.890 113.090 41.290 113.490 ;
        RECT 42.890 113.090 43.290 113.490 ;
        RECT 44.890 113.090 45.290 113.490 ;
        RECT 46.890 113.090 47.290 113.490 ;
        RECT 48.890 113.090 49.290 113.490 ;
        RECT 50.890 113.090 51.290 113.490 ;
        RECT 52.890 113.090 53.290 113.490 ;
        RECT 54.890 113.090 55.290 113.490 ;
        RECT 56.890 113.090 57.290 113.490 ;
        RECT 58.890 113.090 59.290 113.490 ;
        RECT 60.890 113.090 61.290 113.490 ;
        RECT 62.890 113.090 63.290 113.490 ;
        RECT 64.890 113.090 65.290 113.490 ;
        RECT 66.890 113.090 67.290 113.490 ;
        RECT 68.890 113.090 69.290 113.490 ;
        RECT 70.890 113.090 71.290 113.490 ;
        RECT 72.890 113.090 73.290 113.490 ;
        RECT 87.825 113.090 88.225 113.490 ;
        RECT 89.825 113.090 90.225 113.490 ;
        RECT 91.825 113.090 92.225 113.490 ;
        RECT 93.825 113.090 94.225 113.490 ;
        RECT 95.825 113.090 96.225 113.490 ;
        RECT 97.825 113.090 98.225 113.490 ;
        RECT 99.825 113.090 100.225 113.490 ;
        RECT 101.825 113.090 102.225 113.490 ;
        RECT 103.825 113.090 104.225 113.490 ;
        RECT 105.825 113.090 106.225 113.490 ;
        RECT 107.825 113.090 108.225 113.490 ;
        RECT 109.825 113.090 110.225 113.490 ;
        RECT 111.825 113.090 112.225 113.490 ;
        RECT 113.825 113.090 114.225 113.490 ;
        RECT 115.825 113.090 116.225 113.490 ;
        RECT 117.825 113.090 118.225 113.490 ;
        RECT 119.825 113.090 120.225 113.490 ;
        RECT 121.825 113.090 122.225 113.490 ;
        RECT 123.825 113.090 124.225 113.490 ;
        RECT 125.825 113.090 126.225 113.490 ;
        RECT 127.825 113.090 128.225 113.490 ;
        RECT 129.825 113.090 130.225 113.490 ;
        RECT 131.825 113.090 132.225 113.490 ;
        RECT 133.825 113.090 134.225 113.490 ;
        RECT 135.825 113.090 136.225 113.490 ;
        RECT 137.825 113.090 138.225 113.490 ;
        RECT 139.825 113.090 140.225 113.490 ;
        RECT 141.825 113.090 142.225 113.490 ;
        RECT 143.825 113.090 144.225 113.490 ;
        RECT 145.825 113.090 146.225 113.490 ;
        RECT 147.825 113.090 148.225 113.490 ;
        RECT 149.825 113.090 150.225 113.490 ;
        RECT 151.825 113.090 152.225 113.490 ;
        RECT 153.825 113.090 154.225 113.490 ;
        RECT 6.890 112.890 8.540 113.090 ;
        RECT 8.890 112.890 74.540 113.090 ;
        RECT 86.575 112.890 152.225 113.090 ;
        RECT 152.575 112.890 154.225 113.090 ;
        RECT 6.890 112.490 7.290 112.890 ;
        RECT 8.890 112.490 9.290 112.890 ;
        RECT 10.890 112.490 11.290 112.890 ;
        RECT 12.890 112.490 13.290 112.890 ;
        RECT 14.890 112.490 15.290 112.890 ;
        RECT 16.890 112.490 17.290 112.890 ;
        RECT 18.890 112.490 19.290 112.890 ;
        RECT 20.890 112.490 21.290 112.890 ;
        RECT 22.890 112.490 23.290 112.890 ;
        RECT 24.890 112.490 25.290 112.890 ;
        RECT 26.890 112.490 27.290 112.890 ;
        RECT 28.890 112.490 29.290 112.890 ;
        RECT 30.890 112.490 31.290 112.890 ;
        RECT 32.890 112.490 33.290 112.890 ;
        RECT 34.890 112.490 35.290 112.890 ;
        RECT 36.890 112.490 37.290 112.890 ;
        RECT 38.890 112.490 39.290 112.890 ;
        RECT 40.890 112.490 41.290 112.890 ;
        RECT 42.890 112.490 43.290 112.890 ;
        RECT 44.890 112.490 45.290 112.890 ;
        RECT 46.890 112.490 47.290 112.890 ;
        RECT 48.890 112.490 49.290 112.890 ;
        RECT 50.890 112.490 51.290 112.890 ;
        RECT 52.890 112.490 53.290 112.890 ;
        RECT 54.890 112.490 55.290 112.890 ;
        RECT 56.890 112.490 57.290 112.890 ;
        RECT 58.890 112.490 59.290 112.890 ;
        RECT 60.890 112.490 61.290 112.890 ;
        RECT 62.890 112.490 63.290 112.890 ;
        RECT 64.890 112.490 65.290 112.890 ;
        RECT 66.890 112.490 67.290 112.890 ;
        RECT 68.890 112.490 69.290 112.890 ;
        RECT 70.890 112.490 71.290 112.890 ;
        RECT 72.890 112.490 73.290 112.890 ;
        RECT 87.825 112.490 88.225 112.890 ;
        RECT 89.825 112.490 90.225 112.890 ;
        RECT 91.825 112.490 92.225 112.890 ;
        RECT 93.825 112.490 94.225 112.890 ;
        RECT 95.825 112.490 96.225 112.890 ;
        RECT 97.825 112.490 98.225 112.890 ;
        RECT 99.825 112.490 100.225 112.890 ;
        RECT 101.825 112.490 102.225 112.890 ;
        RECT 103.825 112.490 104.225 112.890 ;
        RECT 105.825 112.490 106.225 112.890 ;
        RECT 107.825 112.490 108.225 112.890 ;
        RECT 109.825 112.490 110.225 112.890 ;
        RECT 111.825 112.490 112.225 112.890 ;
        RECT 113.825 112.490 114.225 112.890 ;
        RECT 115.825 112.490 116.225 112.890 ;
        RECT 117.825 112.490 118.225 112.890 ;
        RECT 119.825 112.490 120.225 112.890 ;
        RECT 121.825 112.490 122.225 112.890 ;
        RECT 123.825 112.490 124.225 112.890 ;
        RECT 125.825 112.490 126.225 112.890 ;
        RECT 127.825 112.490 128.225 112.890 ;
        RECT 129.825 112.490 130.225 112.890 ;
        RECT 131.825 112.490 132.225 112.890 ;
        RECT 133.825 112.490 134.225 112.890 ;
        RECT 135.825 112.490 136.225 112.890 ;
        RECT 137.825 112.490 138.225 112.890 ;
        RECT 139.825 112.490 140.225 112.890 ;
        RECT 141.825 112.490 142.225 112.890 ;
        RECT 143.825 112.490 144.225 112.890 ;
        RECT 145.825 112.490 146.225 112.890 ;
        RECT 147.825 112.490 148.225 112.890 ;
        RECT 149.825 112.490 150.225 112.890 ;
        RECT 151.825 112.490 152.225 112.890 ;
        RECT 153.825 112.490 154.225 112.890 ;
        RECT 6.960 111.640 7.220 112.490 ;
        RECT 8.990 111.640 9.190 112.490 ;
        RECT 10.990 111.640 11.190 112.490 ;
        RECT 12.990 111.640 13.190 112.490 ;
        RECT 14.990 111.640 15.190 112.490 ;
        RECT 16.990 111.640 17.190 112.490 ;
        RECT 18.990 111.640 19.190 112.490 ;
        RECT 20.990 111.640 21.190 112.490 ;
        RECT 22.990 111.640 23.190 112.490 ;
        RECT 24.990 111.640 25.190 112.490 ;
        RECT 26.990 111.640 27.190 112.490 ;
        RECT 28.990 111.640 29.190 112.490 ;
        RECT 30.990 111.640 31.190 112.490 ;
        RECT 32.990 111.640 33.190 112.490 ;
        RECT 34.990 111.640 35.190 112.490 ;
        RECT 36.990 111.640 37.190 112.490 ;
        RECT 38.990 111.640 39.190 112.490 ;
        RECT 40.990 111.640 41.190 112.490 ;
        RECT 42.990 111.640 43.190 112.490 ;
        RECT 44.990 111.640 45.190 112.490 ;
        RECT 46.990 111.640 47.190 112.490 ;
        RECT 48.990 111.640 49.190 112.490 ;
        RECT 50.990 111.640 51.190 112.490 ;
        RECT 52.990 111.640 53.190 112.490 ;
        RECT 54.990 111.640 55.190 112.490 ;
        RECT 56.990 111.640 57.190 112.490 ;
        RECT 58.990 111.640 59.190 112.490 ;
        RECT 60.990 111.640 61.190 112.490 ;
        RECT 62.990 111.640 63.190 112.490 ;
        RECT 64.990 111.640 65.190 112.490 ;
        RECT 66.990 111.640 67.190 112.490 ;
        RECT 68.990 111.640 69.190 112.490 ;
        RECT 70.990 111.640 71.190 112.490 ;
        RECT 89.925 111.640 90.125 112.490 ;
        RECT 91.925 111.640 92.125 112.490 ;
        RECT 93.925 111.640 94.125 112.490 ;
        RECT 95.925 111.640 96.125 112.490 ;
        RECT 97.925 111.640 98.125 112.490 ;
        RECT 99.925 111.640 100.125 112.490 ;
        RECT 101.925 111.640 102.125 112.490 ;
        RECT 103.925 111.640 104.125 112.490 ;
        RECT 105.925 111.640 106.125 112.490 ;
        RECT 107.925 111.640 108.125 112.490 ;
        RECT 109.925 111.640 110.125 112.490 ;
        RECT 111.925 111.640 112.125 112.490 ;
        RECT 113.925 111.640 114.125 112.490 ;
        RECT 115.925 111.640 116.125 112.490 ;
        RECT 117.925 111.640 118.125 112.490 ;
        RECT 119.925 111.640 120.125 112.490 ;
        RECT 121.925 111.640 122.125 112.490 ;
        RECT 123.925 111.640 124.125 112.490 ;
        RECT 125.925 111.640 126.125 112.490 ;
        RECT 127.925 111.640 128.125 112.490 ;
        RECT 129.925 111.640 130.125 112.490 ;
        RECT 131.925 111.640 132.125 112.490 ;
        RECT 133.925 111.640 134.125 112.490 ;
        RECT 135.925 111.640 136.125 112.490 ;
        RECT 137.925 111.640 138.125 112.490 ;
        RECT 139.925 111.640 140.125 112.490 ;
        RECT 141.925 111.640 142.125 112.490 ;
        RECT 143.925 111.640 144.125 112.490 ;
        RECT 145.925 111.640 146.125 112.490 ;
        RECT 147.925 111.640 148.125 112.490 ;
        RECT 149.925 111.640 150.125 112.490 ;
        RECT 151.925 111.640 152.125 112.490 ;
        RECT 153.895 111.640 154.155 112.490 ;
        RECT 6.890 111.240 7.290 111.640 ;
        RECT 8.890 111.240 9.290 111.640 ;
        RECT 10.890 111.240 11.290 111.640 ;
        RECT 12.890 111.240 13.290 111.640 ;
        RECT 14.890 111.240 15.290 111.640 ;
        RECT 16.890 111.240 17.290 111.640 ;
        RECT 18.890 111.240 19.290 111.640 ;
        RECT 20.890 111.240 21.290 111.640 ;
        RECT 22.890 111.240 23.290 111.640 ;
        RECT 24.890 111.240 25.290 111.640 ;
        RECT 26.890 111.240 27.290 111.640 ;
        RECT 28.890 111.240 29.290 111.640 ;
        RECT 30.890 111.240 31.290 111.640 ;
        RECT 32.890 111.240 33.290 111.640 ;
        RECT 34.890 111.240 35.290 111.640 ;
        RECT 36.890 111.240 37.290 111.640 ;
        RECT 38.890 111.240 39.290 111.640 ;
        RECT 40.890 111.240 41.290 111.640 ;
        RECT 42.890 111.240 43.290 111.640 ;
        RECT 44.890 111.240 45.290 111.640 ;
        RECT 46.890 111.240 47.290 111.640 ;
        RECT 48.890 111.240 49.290 111.640 ;
        RECT 50.890 111.240 51.290 111.640 ;
        RECT 52.890 111.240 53.290 111.640 ;
        RECT 54.890 111.240 55.290 111.640 ;
        RECT 56.890 111.240 57.290 111.640 ;
        RECT 58.890 111.240 59.290 111.640 ;
        RECT 60.890 111.240 61.290 111.640 ;
        RECT 62.890 111.240 63.290 111.640 ;
        RECT 64.890 111.240 65.290 111.640 ;
        RECT 66.890 111.240 67.290 111.640 ;
        RECT 68.890 111.240 69.290 111.640 ;
        RECT 70.890 111.240 71.290 111.640 ;
        RECT 72.890 111.240 73.290 111.640 ;
        RECT 87.825 111.240 88.225 111.640 ;
        RECT 89.825 111.240 90.225 111.640 ;
        RECT 91.825 111.240 92.225 111.640 ;
        RECT 93.825 111.240 94.225 111.640 ;
        RECT 95.825 111.240 96.225 111.640 ;
        RECT 97.825 111.240 98.225 111.640 ;
        RECT 99.825 111.240 100.225 111.640 ;
        RECT 101.825 111.240 102.225 111.640 ;
        RECT 103.825 111.240 104.225 111.640 ;
        RECT 105.825 111.240 106.225 111.640 ;
        RECT 107.825 111.240 108.225 111.640 ;
        RECT 109.825 111.240 110.225 111.640 ;
        RECT 111.825 111.240 112.225 111.640 ;
        RECT 113.825 111.240 114.225 111.640 ;
        RECT 115.825 111.240 116.225 111.640 ;
        RECT 117.825 111.240 118.225 111.640 ;
        RECT 119.825 111.240 120.225 111.640 ;
        RECT 121.825 111.240 122.225 111.640 ;
        RECT 123.825 111.240 124.225 111.640 ;
        RECT 125.825 111.240 126.225 111.640 ;
        RECT 127.825 111.240 128.225 111.640 ;
        RECT 129.825 111.240 130.225 111.640 ;
        RECT 131.825 111.240 132.225 111.640 ;
        RECT 133.825 111.240 134.225 111.640 ;
        RECT 135.825 111.240 136.225 111.640 ;
        RECT 137.825 111.240 138.225 111.640 ;
        RECT 139.825 111.240 140.225 111.640 ;
        RECT 141.825 111.240 142.225 111.640 ;
        RECT 143.825 111.240 144.225 111.640 ;
        RECT 145.825 111.240 146.225 111.640 ;
        RECT 147.825 111.240 148.225 111.640 ;
        RECT 149.825 111.240 150.225 111.640 ;
        RECT 151.825 111.240 152.225 111.640 ;
        RECT 153.825 111.240 154.225 111.640 ;
        RECT 6.890 111.040 8.540 111.240 ;
        RECT 8.890 111.040 74.540 111.240 ;
        RECT 86.575 111.040 152.225 111.240 ;
        RECT 152.575 111.040 154.225 111.240 ;
        RECT 6.890 110.640 7.290 111.040 ;
        RECT 8.890 110.640 9.290 111.040 ;
        RECT 10.890 110.640 11.290 111.040 ;
        RECT 12.890 110.640 13.290 111.040 ;
        RECT 14.890 110.640 15.290 111.040 ;
        RECT 16.890 110.640 17.290 111.040 ;
        RECT 18.890 110.640 19.290 111.040 ;
        RECT 20.890 110.640 21.290 111.040 ;
        RECT 22.890 110.640 23.290 111.040 ;
        RECT 24.890 110.640 25.290 111.040 ;
        RECT 26.890 110.640 27.290 111.040 ;
        RECT 28.890 110.640 29.290 111.040 ;
        RECT 30.890 110.640 31.290 111.040 ;
        RECT 32.890 110.640 33.290 111.040 ;
        RECT 34.890 110.640 35.290 111.040 ;
        RECT 36.890 110.640 37.290 111.040 ;
        RECT 38.890 110.640 39.290 111.040 ;
        RECT 40.890 110.640 41.290 111.040 ;
        RECT 42.890 110.640 43.290 111.040 ;
        RECT 44.890 110.640 45.290 111.040 ;
        RECT 46.890 110.640 47.290 111.040 ;
        RECT 48.890 110.640 49.290 111.040 ;
        RECT 50.890 110.640 51.290 111.040 ;
        RECT 52.890 110.640 53.290 111.040 ;
        RECT 54.890 110.640 55.290 111.040 ;
        RECT 56.890 110.640 57.290 111.040 ;
        RECT 58.890 110.640 59.290 111.040 ;
        RECT 60.890 110.640 61.290 111.040 ;
        RECT 62.890 110.640 63.290 111.040 ;
        RECT 64.890 110.640 65.290 111.040 ;
        RECT 66.890 110.640 67.290 111.040 ;
        RECT 68.890 110.640 69.290 111.040 ;
        RECT 70.890 110.640 71.290 111.040 ;
        RECT 72.890 110.640 73.290 111.040 ;
        RECT 87.825 110.640 88.225 111.040 ;
        RECT 89.825 110.640 90.225 111.040 ;
        RECT 91.825 110.640 92.225 111.040 ;
        RECT 93.825 110.640 94.225 111.040 ;
        RECT 95.825 110.640 96.225 111.040 ;
        RECT 97.825 110.640 98.225 111.040 ;
        RECT 99.825 110.640 100.225 111.040 ;
        RECT 101.825 110.640 102.225 111.040 ;
        RECT 103.825 110.640 104.225 111.040 ;
        RECT 105.825 110.640 106.225 111.040 ;
        RECT 107.825 110.640 108.225 111.040 ;
        RECT 109.825 110.640 110.225 111.040 ;
        RECT 111.825 110.640 112.225 111.040 ;
        RECT 113.825 110.640 114.225 111.040 ;
        RECT 115.825 110.640 116.225 111.040 ;
        RECT 117.825 110.640 118.225 111.040 ;
        RECT 119.825 110.640 120.225 111.040 ;
        RECT 121.825 110.640 122.225 111.040 ;
        RECT 123.825 110.640 124.225 111.040 ;
        RECT 125.825 110.640 126.225 111.040 ;
        RECT 127.825 110.640 128.225 111.040 ;
        RECT 129.825 110.640 130.225 111.040 ;
        RECT 131.825 110.640 132.225 111.040 ;
        RECT 133.825 110.640 134.225 111.040 ;
        RECT 135.825 110.640 136.225 111.040 ;
        RECT 137.825 110.640 138.225 111.040 ;
        RECT 139.825 110.640 140.225 111.040 ;
        RECT 141.825 110.640 142.225 111.040 ;
        RECT 143.825 110.640 144.225 111.040 ;
        RECT 145.825 110.640 146.225 111.040 ;
        RECT 147.825 110.640 148.225 111.040 ;
        RECT 149.825 110.640 150.225 111.040 ;
        RECT 151.825 110.640 152.225 111.040 ;
        RECT 153.825 110.640 154.225 111.040 ;
        RECT 6.960 109.790 7.220 110.640 ;
        RECT 8.990 109.790 9.190 110.640 ;
        RECT 10.990 109.790 11.190 110.640 ;
        RECT 12.990 109.790 13.190 110.640 ;
        RECT 14.990 109.790 15.190 110.640 ;
        RECT 16.990 109.790 17.190 110.640 ;
        RECT 18.990 109.790 19.190 110.640 ;
        RECT 20.990 109.790 21.190 110.640 ;
        RECT 22.990 109.790 23.190 110.640 ;
        RECT 24.990 109.790 25.190 110.640 ;
        RECT 26.990 109.790 27.190 110.640 ;
        RECT 28.990 109.790 29.190 110.640 ;
        RECT 30.990 109.790 31.190 110.640 ;
        RECT 32.990 109.790 33.190 110.640 ;
        RECT 34.990 109.790 35.190 110.640 ;
        RECT 36.990 109.790 37.190 110.640 ;
        RECT 38.990 109.790 39.190 110.640 ;
        RECT 40.990 109.790 41.190 110.640 ;
        RECT 42.990 109.790 43.190 110.640 ;
        RECT 44.990 109.790 45.190 110.640 ;
        RECT 46.990 109.790 47.190 110.640 ;
        RECT 48.990 109.790 49.190 110.640 ;
        RECT 50.990 109.790 51.190 110.640 ;
        RECT 52.990 109.790 53.190 110.640 ;
        RECT 54.990 109.790 55.190 110.640 ;
        RECT 56.990 109.790 57.190 110.640 ;
        RECT 58.990 109.790 59.190 110.640 ;
        RECT 60.990 109.790 61.190 110.640 ;
        RECT 62.990 109.790 63.190 110.640 ;
        RECT 64.990 109.790 65.190 110.640 ;
        RECT 66.990 109.790 67.190 110.640 ;
        RECT 68.990 109.790 69.190 110.640 ;
        RECT 70.990 109.790 71.190 110.640 ;
        RECT 89.925 109.790 90.125 110.640 ;
        RECT 91.925 109.790 92.125 110.640 ;
        RECT 93.925 109.790 94.125 110.640 ;
        RECT 95.925 109.790 96.125 110.640 ;
        RECT 97.925 109.790 98.125 110.640 ;
        RECT 99.925 109.790 100.125 110.640 ;
        RECT 101.925 109.790 102.125 110.640 ;
        RECT 103.925 109.790 104.125 110.640 ;
        RECT 105.925 109.790 106.125 110.640 ;
        RECT 107.925 109.790 108.125 110.640 ;
        RECT 109.925 109.790 110.125 110.640 ;
        RECT 111.925 109.790 112.125 110.640 ;
        RECT 113.925 109.790 114.125 110.640 ;
        RECT 115.925 109.790 116.125 110.640 ;
        RECT 117.925 109.790 118.125 110.640 ;
        RECT 119.925 109.790 120.125 110.640 ;
        RECT 121.925 109.790 122.125 110.640 ;
        RECT 123.925 109.790 124.125 110.640 ;
        RECT 125.925 109.790 126.125 110.640 ;
        RECT 127.925 109.790 128.125 110.640 ;
        RECT 129.925 109.790 130.125 110.640 ;
        RECT 131.925 109.790 132.125 110.640 ;
        RECT 133.925 109.790 134.125 110.640 ;
        RECT 135.925 109.790 136.125 110.640 ;
        RECT 137.925 109.790 138.125 110.640 ;
        RECT 139.925 109.790 140.125 110.640 ;
        RECT 141.925 109.790 142.125 110.640 ;
        RECT 143.925 109.790 144.125 110.640 ;
        RECT 145.925 109.790 146.125 110.640 ;
        RECT 147.925 109.790 148.125 110.640 ;
        RECT 149.925 109.790 150.125 110.640 ;
        RECT 151.925 109.790 152.125 110.640 ;
        RECT 153.895 109.790 154.155 110.640 ;
        RECT 6.890 109.390 7.290 109.790 ;
        RECT 8.890 109.390 9.290 109.790 ;
        RECT 10.890 109.390 11.290 109.790 ;
        RECT 12.890 109.390 13.290 109.790 ;
        RECT 14.890 109.390 15.290 109.790 ;
        RECT 16.890 109.390 17.290 109.790 ;
        RECT 18.890 109.390 19.290 109.790 ;
        RECT 20.890 109.390 21.290 109.790 ;
        RECT 22.890 109.390 23.290 109.790 ;
        RECT 24.890 109.390 25.290 109.790 ;
        RECT 26.890 109.390 27.290 109.790 ;
        RECT 28.890 109.390 29.290 109.790 ;
        RECT 30.890 109.390 31.290 109.790 ;
        RECT 32.890 109.390 33.290 109.790 ;
        RECT 34.890 109.390 35.290 109.790 ;
        RECT 36.890 109.390 37.290 109.790 ;
        RECT 38.890 109.390 39.290 109.790 ;
        RECT 40.890 109.390 41.290 109.790 ;
        RECT 42.890 109.390 43.290 109.790 ;
        RECT 44.890 109.390 45.290 109.790 ;
        RECT 46.890 109.390 47.290 109.790 ;
        RECT 48.890 109.390 49.290 109.790 ;
        RECT 50.890 109.390 51.290 109.790 ;
        RECT 52.890 109.390 53.290 109.790 ;
        RECT 54.890 109.390 55.290 109.790 ;
        RECT 56.890 109.390 57.290 109.790 ;
        RECT 58.890 109.390 59.290 109.790 ;
        RECT 60.890 109.390 61.290 109.790 ;
        RECT 62.890 109.390 63.290 109.790 ;
        RECT 64.890 109.390 65.290 109.790 ;
        RECT 66.890 109.390 67.290 109.790 ;
        RECT 68.890 109.390 69.290 109.790 ;
        RECT 70.890 109.390 71.290 109.790 ;
        RECT 72.890 109.390 73.290 109.790 ;
        RECT 87.825 109.390 88.225 109.790 ;
        RECT 89.825 109.390 90.225 109.790 ;
        RECT 91.825 109.390 92.225 109.790 ;
        RECT 93.825 109.390 94.225 109.790 ;
        RECT 95.825 109.390 96.225 109.790 ;
        RECT 97.825 109.390 98.225 109.790 ;
        RECT 99.825 109.390 100.225 109.790 ;
        RECT 101.825 109.390 102.225 109.790 ;
        RECT 103.825 109.390 104.225 109.790 ;
        RECT 105.825 109.390 106.225 109.790 ;
        RECT 107.825 109.390 108.225 109.790 ;
        RECT 109.825 109.390 110.225 109.790 ;
        RECT 111.825 109.390 112.225 109.790 ;
        RECT 113.825 109.390 114.225 109.790 ;
        RECT 115.825 109.390 116.225 109.790 ;
        RECT 117.825 109.390 118.225 109.790 ;
        RECT 119.825 109.390 120.225 109.790 ;
        RECT 121.825 109.390 122.225 109.790 ;
        RECT 123.825 109.390 124.225 109.790 ;
        RECT 125.825 109.390 126.225 109.790 ;
        RECT 127.825 109.390 128.225 109.790 ;
        RECT 129.825 109.390 130.225 109.790 ;
        RECT 131.825 109.390 132.225 109.790 ;
        RECT 133.825 109.390 134.225 109.790 ;
        RECT 135.825 109.390 136.225 109.790 ;
        RECT 137.825 109.390 138.225 109.790 ;
        RECT 139.825 109.390 140.225 109.790 ;
        RECT 141.825 109.390 142.225 109.790 ;
        RECT 143.825 109.390 144.225 109.790 ;
        RECT 145.825 109.390 146.225 109.790 ;
        RECT 147.825 109.390 148.225 109.790 ;
        RECT 149.825 109.390 150.225 109.790 ;
        RECT 151.825 109.390 152.225 109.790 ;
        RECT 153.825 109.390 154.225 109.790 ;
        RECT 6.890 109.190 8.540 109.390 ;
        RECT 8.890 109.190 74.540 109.390 ;
        RECT 86.575 109.190 152.225 109.390 ;
        RECT 152.575 109.190 154.225 109.390 ;
        RECT 6.890 108.790 7.290 109.190 ;
        RECT 8.890 108.790 9.290 109.190 ;
        RECT 10.890 108.790 11.290 109.190 ;
        RECT 12.890 108.790 13.290 109.190 ;
        RECT 14.890 108.790 15.290 109.190 ;
        RECT 16.890 108.790 17.290 109.190 ;
        RECT 18.890 108.790 19.290 109.190 ;
        RECT 20.890 108.790 21.290 109.190 ;
        RECT 22.890 108.790 23.290 109.190 ;
        RECT 24.890 108.790 25.290 109.190 ;
        RECT 26.890 108.790 27.290 109.190 ;
        RECT 28.890 108.790 29.290 109.190 ;
        RECT 30.890 108.790 31.290 109.190 ;
        RECT 32.890 108.790 33.290 109.190 ;
        RECT 34.890 108.790 35.290 109.190 ;
        RECT 36.890 108.790 37.290 109.190 ;
        RECT 38.890 108.790 39.290 109.190 ;
        RECT 40.890 108.790 41.290 109.190 ;
        RECT 42.890 108.790 43.290 109.190 ;
        RECT 44.890 108.790 45.290 109.190 ;
        RECT 46.890 108.790 47.290 109.190 ;
        RECT 48.890 108.790 49.290 109.190 ;
        RECT 50.890 108.790 51.290 109.190 ;
        RECT 52.890 108.790 53.290 109.190 ;
        RECT 54.890 108.790 55.290 109.190 ;
        RECT 56.890 108.790 57.290 109.190 ;
        RECT 58.890 108.790 59.290 109.190 ;
        RECT 60.890 108.790 61.290 109.190 ;
        RECT 62.890 108.790 63.290 109.190 ;
        RECT 64.890 108.790 65.290 109.190 ;
        RECT 66.890 108.790 67.290 109.190 ;
        RECT 68.890 108.790 69.290 109.190 ;
        RECT 70.890 108.790 71.290 109.190 ;
        RECT 72.890 108.790 73.290 109.190 ;
        RECT 87.825 108.790 88.225 109.190 ;
        RECT 89.825 108.790 90.225 109.190 ;
        RECT 91.825 108.790 92.225 109.190 ;
        RECT 93.825 108.790 94.225 109.190 ;
        RECT 95.825 108.790 96.225 109.190 ;
        RECT 97.825 108.790 98.225 109.190 ;
        RECT 99.825 108.790 100.225 109.190 ;
        RECT 101.825 108.790 102.225 109.190 ;
        RECT 103.825 108.790 104.225 109.190 ;
        RECT 105.825 108.790 106.225 109.190 ;
        RECT 107.825 108.790 108.225 109.190 ;
        RECT 109.825 108.790 110.225 109.190 ;
        RECT 111.825 108.790 112.225 109.190 ;
        RECT 113.825 108.790 114.225 109.190 ;
        RECT 115.825 108.790 116.225 109.190 ;
        RECT 117.825 108.790 118.225 109.190 ;
        RECT 119.825 108.790 120.225 109.190 ;
        RECT 121.825 108.790 122.225 109.190 ;
        RECT 123.825 108.790 124.225 109.190 ;
        RECT 125.825 108.790 126.225 109.190 ;
        RECT 127.825 108.790 128.225 109.190 ;
        RECT 129.825 108.790 130.225 109.190 ;
        RECT 131.825 108.790 132.225 109.190 ;
        RECT 133.825 108.790 134.225 109.190 ;
        RECT 135.825 108.790 136.225 109.190 ;
        RECT 137.825 108.790 138.225 109.190 ;
        RECT 139.825 108.790 140.225 109.190 ;
        RECT 141.825 108.790 142.225 109.190 ;
        RECT 143.825 108.790 144.225 109.190 ;
        RECT 145.825 108.790 146.225 109.190 ;
        RECT 147.825 108.790 148.225 109.190 ;
        RECT 149.825 108.790 150.225 109.190 ;
        RECT 151.825 108.790 152.225 109.190 ;
        RECT 153.825 108.790 154.225 109.190 ;
        RECT 6.960 107.940 7.220 108.790 ;
        RECT 8.990 107.940 9.190 108.790 ;
        RECT 10.990 107.940 11.190 108.790 ;
        RECT 12.990 107.940 13.190 108.790 ;
        RECT 14.990 107.940 15.190 108.790 ;
        RECT 16.990 107.940 17.190 108.790 ;
        RECT 18.990 107.940 19.190 108.790 ;
        RECT 20.990 107.940 21.190 108.790 ;
        RECT 22.990 107.940 23.190 108.790 ;
        RECT 24.990 107.940 25.190 108.790 ;
        RECT 26.990 107.940 27.190 108.790 ;
        RECT 28.990 107.940 29.190 108.790 ;
        RECT 30.990 107.940 31.190 108.790 ;
        RECT 32.990 107.940 33.190 108.790 ;
        RECT 34.990 107.940 35.190 108.790 ;
        RECT 36.990 107.940 37.190 108.790 ;
        RECT 38.990 107.940 39.190 108.790 ;
        RECT 40.990 107.940 41.190 108.790 ;
        RECT 42.990 107.940 43.190 108.790 ;
        RECT 44.990 107.940 45.190 108.790 ;
        RECT 46.990 107.940 47.190 108.790 ;
        RECT 48.990 107.940 49.190 108.790 ;
        RECT 50.990 107.940 51.190 108.790 ;
        RECT 52.990 107.940 53.190 108.790 ;
        RECT 54.990 107.940 55.190 108.790 ;
        RECT 56.990 107.940 57.190 108.790 ;
        RECT 58.990 107.940 59.190 108.790 ;
        RECT 60.990 107.940 61.190 108.790 ;
        RECT 62.990 107.940 63.190 108.790 ;
        RECT 64.990 107.940 65.190 108.790 ;
        RECT 66.990 107.940 67.190 108.790 ;
        RECT 68.990 107.940 69.190 108.790 ;
        RECT 70.990 107.940 71.190 108.790 ;
        RECT 89.925 107.940 90.125 108.790 ;
        RECT 91.925 107.940 92.125 108.790 ;
        RECT 93.925 107.940 94.125 108.790 ;
        RECT 95.925 107.940 96.125 108.790 ;
        RECT 97.925 107.940 98.125 108.790 ;
        RECT 99.925 107.940 100.125 108.790 ;
        RECT 101.925 107.940 102.125 108.790 ;
        RECT 103.925 107.940 104.125 108.790 ;
        RECT 105.925 107.940 106.125 108.790 ;
        RECT 107.925 107.940 108.125 108.790 ;
        RECT 109.925 107.940 110.125 108.790 ;
        RECT 111.925 107.940 112.125 108.790 ;
        RECT 113.925 107.940 114.125 108.790 ;
        RECT 115.925 107.940 116.125 108.790 ;
        RECT 117.925 107.940 118.125 108.790 ;
        RECT 119.925 107.940 120.125 108.790 ;
        RECT 121.925 107.940 122.125 108.790 ;
        RECT 123.925 107.940 124.125 108.790 ;
        RECT 125.925 107.940 126.125 108.790 ;
        RECT 127.925 107.940 128.125 108.790 ;
        RECT 129.925 107.940 130.125 108.790 ;
        RECT 131.925 107.940 132.125 108.790 ;
        RECT 133.925 107.940 134.125 108.790 ;
        RECT 135.925 107.940 136.125 108.790 ;
        RECT 137.925 107.940 138.125 108.790 ;
        RECT 139.925 107.940 140.125 108.790 ;
        RECT 141.925 107.940 142.125 108.790 ;
        RECT 143.925 107.940 144.125 108.790 ;
        RECT 145.925 107.940 146.125 108.790 ;
        RECT 147.925 107.940 148.125 108.790 ;
        RECT 149.925 107.940 150.125 108.790 ;
        RECT 151.925 107.940 152.125 108.790 ;
        RECT 153.895 107.940 154.155 108.790 ;
        RECT 6.890 107.540 7.290 107.940 ;
        RECT 8.890 107.540 9.290 107.940 ;
        RECT 10.890 107.540 11.290 107.940 ;
        RECT 12.890 107.540 13.290 107.940 ;
        RECT 14.890 107.540 15.290 107.940 ;
        RECT 16.890 107.540 17.290 107.940 ;
        RECT 18.890 107.540 19.290 107.940 ;
        RECT 20.890 107.540 21.290 107.940 ;
        RECT 22.890 107.540 23.290 107.940 ;
        RECT 24.890 107.540 25.290 107.940 ;
        RECT 26.890 107.540 27.290 107.940 ;
        RECT 28.890 107.540 29.290 107.940 ;
        RECT 30.890 107.540 31.290 107.940 ;
        RECT 32.890 107.540 33.290 107.940 ;
        RECT 34.890 107.540 35.290 107.940 ;
        RECT 36.890 107.540 37.290 107.940 ;
        RECT 38.890 107.540 39.290 107.940 ;
        RECT 40.890 107.540 41.290 107.940 ;
        RECT 42.890 107.540 43.290 107.940 ;
        RECT 44.890 107.540 45.290 107.940 ;
        RECT 46.890 107.540 47.290 107.940 ;
        RECT 48.890 107.540 49.290 107.940 ;
        RECT 50.890 107.540 51.290 107.940 ;
        RECT 52.890 107.540 53.290 107.940 ;
        RECT 54.890 107.540 55.290 107.940 ;
        RECT 56.890 107.540 57.290 107.940 ;
        RECT 58.890 107.540 59.290 107.940 ;
        RECT 60.890 107.540 61.290 107.940 ;
        RECT 62.890 107.540 63.290 107.940 ;
        RECT 64.890 107.540 65.290 107.940 ;
        RECT 66.890 107.540 67.290 107.940 ;
        RECT 68.890 107.540 69.290 107.940 ;
        RECT 70.890 107.540 71.290 107.940 ;
        RECT 72.890 107.540 73.290 107.940 ;
        RECT 87.825 107.540 88.225 107.940 ;
        RECT 89.825 107.540 90.225 107.940 ;
        RECT 91.825 107.540 92.225 107.940 ;
        RECT 93.825 107.540 94.225 107.940 ;
        RECT 95.825 107.540 96.225 107.940 ;
        RECT 97.825 107.540 98.225 107.940 ;
        RECT 99.825 107.540 100.225 107.940 ;
        RECT 101.825 107.540 102.225 107.940 ;
        RECT 103.825 107.540 104.225 107.940 ;
        RECT 105.825 107.540 106.225 107.940 ;
        RECT 107.825 107.540 108.225 107.940 ;
        RECT 109.825 107.540 110.225 107.940 ;
        RECT 111.825 107.540 112.225 107.940 ;
        RECT 113.825 107.540 114.225 107.940 ;
        RECT 115.825 107.540 116.225 107.940 ;
        RECT 117.825 107.540 118.225 107.940 ;
        RECT 119.825 107.540 120.225 107.940 ;
        RECT 121.825 107.540 122.225 107.940 ;
        RECT 123.825 107.540 124.225 107.940 ;
        RECT 125.825 107.540 126.225 107.940 ;
        RECT 127.825 107.540 128.225 107.940 ;
        RECT 129.825 107.540 130.225 107.940 ;
        RECT 131.825 107.540 132.225 107.940 ;
        RECT 133.825 107.540 134.225 107.940 ;
        RECT 135.825 107.540 136.225 107.940 ;
        RECT 137.825 107.540 138.225 107.940 ;
        RECT 139.825 107.540 140.225 107.940 ;
        RECT 141.825 107.540 142.225 107.940 ;
        RECT 143.825 107.540 144.225 107.940 ;
        RECT 145.825 107.540 146.225 107.940 ;
        RECT 147.825 107.540 148.225 107.940 ;
        RECT 149.825 107.540 150.225 107.940 ;
        RECT 151.825 107.540 152.225 107.940 ;
        RECT 153.825 107.540 154.225 107.940 ;
        RECT 6.890 107.340 8.540 107.540 ;
        RECT 8.890 107.340 74.540 107.540 ;
        RECT 86.575 107.340 152.225 107.540 ;
        RECT 152.575 107.340 154.225 107.540 ;
        RECT 6.890 106.940 7.290 107.340 ;
        RECT 8.890 106.940 9.290 107.340 ;
        RECT 10.890 106.940 11.290 107.340 ;
        RECT 12.890 106.940 13.290 107.340 ;
        RECT 14.890 106.940 15.290 107.340 ;
        RECT 16.890 106.940 17.290 107.340 ;
        RECT 18.890 106.940 19.290 107.340 ;
        RECT 20.890 106.940 21.290 107.340 ;
        RECT 22.890 106.940 23.290 107.340 ;
        RECT 24.890 106.940 25.290 107.340 ;
        RECT 26.890 106.940 27.290 107.340 ;
        RECT 28.890 106.940 29.290 107.340 ;
        RECT 30.890 106.940 31.290 107.340 ;
        RECT 32.890 106.940 33.290 107.340 ;
        RECT 34.890 106.940 35.290 107.340 ;
        RECT 36.890 106.940 37.290 107.340 ;
        RECT 38.890 106.940 39.290 107.340 ;
        RECT 40.890 106.940 41.290 107.340 ;
        RECT 42.890 106.940 43.290 107.340 ;
        RECT 44.890 106.940 45.290 107.340 ;
        RECT 46.890 106.940 47.290 107.340 ;
        RECT 48.890 106.940 49.290 107.340 ;
        RECT 50.890 106.940 51.290 107.340 ;
        RECT 52.890 106.940 53.290 107.340 ;
        RECT 54.890 106.940 55.290 107.340 ;
        RECT 56.890 106.940 57.290 107.340 ;
        RECT 58.890 106.940 59.290 107.340 ;
        RECT 60.890 106.940 61.290 107.340 ;
        RECT 62.890 106.940 63.290 107.340 ;
        RECT 64.890 106.940 65.290 107.340 ;
        RECT 66.890 106.940 67.290 107.340 ;
        RECT 68.890 106.940 69.290 107.340 ;
        RECT 70.890 106.940 71.290 107.340 ;
        RECT 72.890 106.940 73.290 107.340 ;
        RECT 87.825 106.940 88.225 107.340 ;
        RECT 89.825 106.940 90.225 107.340 ;
        RECT 91.825 106.940 92.225 107.340 ;
        RECT 93.825 106.940 94.225 107.340 ;
        RECT 95.825 106.940 96.225 107.340 ;
        RECT 97.825 106.940 98.225 107.340 ;
        RECT 99.825 106.940 100.225 107.340 ;
        RECT 101.825 106.940 102.225 107.340 ;
        RECT 103.825 106.940 104.225 107.340 ;
        RECT 105.825 106.940 106.225 107.340 ;
        RECT 107.825 106.940 108.225 107.340 ;
        RECT 109.825 106.940 110.225 107.340 ;
        RECT 111.825 106.940 112.225 107.340 ;
        RECT 113.825 106.940 114.225 107.340 ;
        RECT 115.825 106.940 116.225 107.340 ;
        RECT 117.825 106.940 118.225 107.340 ;
        RECT 119.825 106.940 120.225 107.340 ;
        RECT 121.825 106.940 122.225 107.340 ;
        RECT 123.825 106.940 124.225 107.340 ;
        RECT 125.825 106.940 126.225 107.340 ;
        RECT 127.825 106.940 128.225 107.340 ;
        RECT 129.825 106.940 130.225 107.340 ;
        RECT 131.825 106.940 132.225 107.340 ;
        RECT 133.825 106.940 134.225 107.340 ;
        RECT 135.825 106.940 136.225 107.340 ;
        RECT 137.825 106.940 138.225 107.340 ;
        RECT 139.825 106.940 140.225 107.340 ;
        RECT 141.825 106.940 142.225 107.340 ;
        RECT 143.825 106.940 144.225 107.340 ;
        RECT 145.825 106.940 146.225 107.340 ;
        RECT 147.825 106.940 148.225 107.340 ;
        RECT 149.825 106.940 150.225 107.340 ;
        RECT 151.825 106.940 152.225 107.340 ;
        RECT 153.825 106.940 154.225 107.340 ;
        RECT 6.960 106.090 7.220 106.940 ;
        RECT 8.990 106.090 9.190 106.940 ;
        RECT 10.990 106.090 11.190 106.940 ;
        RECT 12.990 106.090 13.190 106.940 ;
        RECT 14.990 106.090 15.190 106.940 ;
        RECT 16.990 106.090 17.190 106.940 ;
        RECT 18.990 106.090 19.190 106.940 ;
        RECT 20.990 106.090 21.190 106.940 ;
        RECT 22.990 106.090 23.190 106.940 ;
        RECT 24.990 106.090 25.190 106.940 ;
        RECT 26.990 106.090 27.190 106.940 ;
        RECT 28.990 106.090 29.190 106.940 ;
        RECT 30.990 106.090 31.190 106.940 ;
        RECT 32.990 106.090 33.190 106.940 ;
        RECT 34.990 106.090 35.190 106.940 ;
        RECT 36.990 106.090 37.190 106.940 ;
        RECT 38.990 106.090 39.190 106.940 ;
        RECT 40.990 106.090 41.190 106.940 ;
        RECT 42.990 106.090 43.190 106.940 ;
        RECT 44.990 106.090 45.190 106.940 ;
        RECT 46.990 106.090 47.190 106.940 ;
        RECT 48.990 106.090 49.190 106.940 ;
        RECT 50.990 106.090 51.190 106.940 ;
        RECT 52.990 106.090 53.190 106.940 ;
        RECT 54.990 106.090 55.190 106.940 ;
        RECT 56.990 106.090 57.190 106.940 ;
        RECT 58.990 106.090 59.190 106.940 ;
        RECT 60.990 106.090 61.190 106.940 ;
        RECT 62.990 106.090 63.190 106.940 ;
        RECT 64.990 106.090 65.190 106.940 ;
        RECT 66.990 106.090 67.190 106.940 ;
        RECT 68.990 106.090 69.190 106.940 ;
        RECT 70.990 106.090 71.190 106.940 ;
        RECT 89.925 106.090 90.125 106.940 ;
        RECT 91.925 106.090 92.125 106.940 ;
        RECT 93.925 106.090 94.125 106.940 ;
        RECT 95.925 106.090 96.125 106.940 ;
        RECT 97.925 106.090 98.125 106.940 ;
        RECT 99.925 106.090 100.125 106.940 ;
        RECT 101.925 106.090 102.125 106.940 ;
        RECT 103.925 106.090 104.125 106.940 ;
        RECT 105.925 106.090 106.125 106.940 ;
        RECT 107.925 106.090 108.125 106.940 ;
        RECT 109.925 106.090 110.125 106.940 ;
        RECT 111.925 106.090 112.125 106.940 ;
        RECT 113.925 106.090 114.125 106.940 ;
        RECT 115.925 106.090 116.125 106.940 ;
        RECT 117.925 106.090 118.125 106.940 ;
        RECT 119.925 106.090 120.125 106.940 ;
        RECT 121.925 106.090 122.125 106.940 ;
        RECT 123.925 106.090 124.125 106.940 ;
        RECT 125.925 106.090 126.125 106.940 ;
        RECT 127.925 106.090 128.125 106.940 ;
        RECT 129.925 106.090 130.125 106.940 ;
        RECT 131.925 106.090 132.125 106.940 ;
        RECT 133.925 106.090 134.125 106.940 ;
        RECT 135.925 106.090 136.125 106.940 ;
        RECT 137.925 106.090 138.125 106.940 ;
        RECT 139.925 106.090 140.125 106.940 ;
        RECT 141.925 106.090 142.125 106.940 ;
        RECT 143.925 106.090 144.125 106.940 ;
        RECT 145.925 106.090 146.125 106.940 ;
        RECT 147.925 106.090 148.125 106.940 ;
        RECT 149.925 106.090 150.125 106.940 ;
        RECT 151.925 106.090 152.125 106.940 ;
        RECT 153.895 106.090 154.155 106.940 ;
        RECT 6.890 105.690 7.290 106.090 ;
        RECT 8.890 105.690 9.290 106.090 ;
        RECT 10.890 105.690 11.290 106.090 ;
        RECT 12.890 105.690 13.290 106.090 ;
        RECT 14.890 105.690 15.290 106.090 ;
        RECT 16.890 105.690 17.290 106.090 ;
        RECT 18.890 105.690 19.290 106.090 ;
        RECT 20.890 105.690 21.290 106.090 ;
        RECT 22.890 105.690 23.290 106.090 ;
        RECT 24.890 105.690 25.290 106.090 ;
        RECT 26.890 105.690 27.290 106.090 ;
        RECT 28.890 105.690 29.290 106.090 ;
        RECT 30.890 105.690 31.290 106.090 ;
        RECT 32.890 105.690 33.290 106.090 ;
        RECT 34.890 105.690 35.290 106.090 ;
        RECT 36.890 105.690 37.290 106.090 ;
        RECT 38.890 105.690 39.290 106.090 ;
        RECT 40.890 105.690 41.290 106.090 ;
        RECT 42.890 105.690 43.290 106.090 ;
        RECT 44.890 105.690 45.290 106.090 ;
        RECT 46.890 105.690 47.290 106.090 ;
        RECT 48.890 105.690 49.290 106.090 ;
        RECT 50.890 105.690 51.290 106.090 ;
        RECT 52.890 105.690 53.290 106.090 ;
        RECT 54.890 105.690 55.290 106.090 ;
        RECT 56.890 105.690 57.290 106.090 ;
        RECT 58.890 105.690 59.290 106.090 ;
        RECT 60.890 105.690 61.290 106.090 ;
        RECT 62.890 105.690 63.290 106.090 ;
        RECT 64.890 105.690 65.290 106.090 ;
        RECT 66.890 105.690 67.290 106.090 ;
        RECT 68.890 105.690 69.290 106.090 ;
        RECT 70.890 105.690 71.290 106.090 ;
        RECT 72.890 105.690 73.290 106.090 ;
        RECT 87.825 105.690 88.225 106.090 ;
        RECT 89.825 105.690 90.225 106.090 ;
        RECT 91.825 105.690 92.225 106.090 ;
        RECT 93.825 105.690 94.225 106.090 ;
        RECT 95.825 105.690 96.225 106.090 ;
        RECT 97.825 105.690 98.225 106.090 ;
        RECT 99.825 105.690 100.225 106.090 ;
        RECT 101.825 105.690 102.225 106.090 ;
        RECT 103.825 105.690 104.225 106.090 ;
        RECT 105.825 105.690 106.225 106.090 ;
        RECT 107.825 105.690 108.225 106.090 ;
        RECT 109.825 105.690 110.225 106.090 ;
        RECT 111.825 105.690 112.225 106.090 ;
        RECT 113.825 105.690 114.225 106.090 ;
        RECT 115.825 105.690 116.225 106.090 ;
        RECT 117.825 105.690 118.225 106.090 ;
        RECT 119.825 105.690 120.225 106.090 ;
        RECT 121.825 105.690 122.225 106.090 ;
        RECT 123.825 105.690 124.225 106.090 ;
        RECT 125.825 105.690 126.225 106.090 ;
        RECT 127.825 105.690 128.225 106.090 ;
        RECT 129.825 105.690 130.225 106.090 ;
        RECT 131.825 105.690 132.225 106.090 ;
        RECT 133.825 105.690 134.225 106.090 ;
        RECT 135.825 105.690 136.225 106.090 ;
        RECT 137.825 105.690 138.225 106.090 ;
        RECT 139.825 105.690 140.225 106.090 ;
        RECT 141.825 105.690 142.225 106.090 ;
        RECT 143.825 105.690 144.225 106.090 ;
        RECT 145.825 105.690 146.225 106.090 ;
        RECT 147.825 105.690 148.225 106.090 ;
        RECT 149.825 105.690 150.225 106.090 ;
        RECT 151.825 105.690 152.225 106.090 ;
        RECT 153.825 105.690 154.225 106.090 ;
        RECT 6.890 105.490 8.540 105.690 ;
        RECT 8.890 105.490 74.540 105.690 ;
        RECT 86.575 105.490 152.225 105.690 ;
        RECT 152.575 105.490 154.225 105.690 ;
        RECT 6.890 105.090 7.290 105.490 ;
        RECT 8.890 105.090 9.290 105.490 ;
        RECT 10.890 105.090 11.290 105.490 ;
        RECT 12.890 105.090 13.290 105.490 ;
        RECT 14.890 105.090 15.290 105.490 ;
        RECT 16.890 105.090 17.290 105.490 ;
        RECT 18.890 105.090 19.290 105.490 ;
        RECT 20.890 105.090 21.290 105.490 ;
        RECT 22.890 105.090 23.290 105.490 ;
        RECT 24.890 105.090 25.290 105.490 ;
        RECT 26.890 105.090 27.290 105.490 ;
        RECT 28.890 105.090 29.290 105.490 ;
        RECT 30.890 105.090 31.290 105.490 ;
        RECT 32.890 105.090 33.290 105.490 ;
        RECT 34.890 105.090 35.290 105.490 ;
        RECT 36.890 105.090 37.290 105.490 ;
        RECT 38.890 105.090 39.290 105.490 ;
        RECT 40.890 105.090 41.290 105.490 ;
        RECT 42.890 105.090 43.290 105.490 ;
        RECT 44.890 105.090 45.290 105.490 ;
        RECT 46.890 105.090 47.290 105.490 ;
        RECT 48.890 105.090 49.290 105.490 ;
        RECT 50.890 105.090 51.290 105.490 ;
        RECT 52.890 105.090 53.290 105.490 ;
        RECT 54.890 105.090 55.290 105.490 ;
        RECT 56.890 105.090 57.290 105.490 ;
        RECT 58.890 105.090 59.290 105.490 ;
        RECT 60.890 105.090 61.290 105.490 ;
        RECT 62.890 105.090 63.290 105.490 ;
        RECT 64.890 105.090 65.290 105.490 ;
        RECT 66.890 105.090 67.290 105.490 ;
        RECT 68.890 105.090 69.290 105.490 ;
        RECT 70.890 105.090 71.290 105.490 ;
        RECT 72.890 105.090 73.290 105.490 ;
        RECT 87.825 105.090 88.225 105.490 ;
        RECT 89.825 105.090 90.225 105.490 ;
        RECT 91.825 105.090 92.225 105.490 ;
        RECT 93.825 105.090 94.225 105.490 ;
        RECT 95.825 105.090 96.225 105.490 ;
        RECT 97.825 105.090 98.225 105.490 ;
        RECT 99.825 105.090 100.225 105.490 ;
        RECT 101.825 105.090 102.225 105.490 ;
        RECT 103.825 105.090 104.225 105.490 ;
        RECT 105.825 105.090 106.225 105.490 ;
        RECT 107.825 105.090 108.225 105.490 ;
        RECT 109.825 105.090 110.225 105.490 ;
        RECT 111.825 105.090 112.225 105.490 ;
        RECT 113.825 105.090 114.225 105.490 ;
        RECT 115.825 105.090 116.225 105.490 ;
        RECT 117.825 105.090 118.225 105.490 ;
        RECT 119.825 105.090 120.225 105.490 ;
        RECT 121.825 105.090 122.225 105.490 ;
        RECT 123.825 105.090 124.225 105.490 ;
        RECT 125.825 105.090 126.225 105.490 ;
        RECT 127.825 105.090 128.225 105.490 ;
        RECT 129.825 105.090 130.225 105.490 ;
        RECT 131.825 105.090 132.225 105.490 ;
        RECT 133.825 105.090 134.225 105.490 ;
        RECT 135.825 105.090 136.225 105.490 ;
        RECT 137.825 105.090 138.225 105.490 ;
        RECT 139.825 105.090 140.225 105.490 ;
        RECT 141.825 105.090 142.225 105.490 ;
        RECT 143.825 105.090 144.225 105.490 ;
        RECT 145.825 105.090 146.225 105.490 ;
        RECT 147.825 105.090 148.225 105.490 ;
        RECT 149.825 105.090 150.225 105.490 ;
        RECT 151.825 105.090 152.225 105.490 ;
        RECT 153.825 105.090 154.225 105.490 ;
        RECT 6.960 104.240 7.220 105.090 ;
        RECT 8.990 104.240 9.190 105.090 ;
        RECT 10.990 104.240 11.190 105.090 ;
        RECT 12.990 104.240 13.190 105.090 ;
        RECT 14.990 104.240 15.190 105.090 ;
        RECT 16.990 104.240 17.190 105.090 ;
        RECT 18.990 104.240 19.190 105.090 ;
        RECT 20.990 104.240 21.190 105.090 ;
        RECT 22.990 104.240 23.190 105.090 ;
        RECT 137.925 104.240 138.125 105.090 ;
        RECT 139.925 104.240 140.125 105.090 ;
        RECT 141.925 104.240 142.125 105.090 ;
        RECT 143.925 104.240 144.125 105.090 ;
        RECT 145.925 104.240 146.125 105.090 ;
        RECT 147.925 104.240 148.125 105.090 ;
        RECT 149.925 104.240 150.125 105.090 ;
        RECT 151.925 104.240 152.125 105.090 ;
        RECT 153.895 104.240 154.155 105.090 ;
        RECT 6.890 103.840 7.290 104.240 ;
        RECT 8.890 103.840 9.290 104.240 ;
        RECT 10.890 103.840 11.290 104.240 ;
        RECT 12.890 103.840 13.290 104.240 ;
        RECT 14.890 103.840 15.290 104.240 ;
        RECT 16.890 103.840 17.290 104.240 ;
        RECT 18.890 103.840 19.290 104.240 ;
        RECT 20.890 103.840 21.290 104.240 ;
        RECT 22.890 103.840 23.290 104.240 ;
        RECT 24.890 103.840 25.290 104.240 ;
        RECT 26.890 103.840 27.290 104.240 ;
        RECT 28.890 103.840 29.290 104.240 ;
        RECT 30.890 103.840 31.290 104.240 ;
        RECT 32.890 103.840 33.290 104.240 ;
        RECT 34.890 103.840 35.290 104.240 ;
        RECT 36.890 103.840 37.290 104.240 ;
        RECT 38.890 103.840 39.290 104.240 ;
        RECT 40.890 103.840 41.290 104.240 ;
        RECT 42.890 103.840 43.290 104.240 ;
        RECT 44.890 103.840 45.290 104.240 ;
        RECT 46.890 103.840 47.290 104.240 ;
        RECT 48.890 103.840 49.290 104.240 ;
        RECT 50.890 103.840 51.290 104.240 ;
        RECT 52.890 103.840 53.290 104.240 ;
        RECT 54.890 103.840 55.290 104.240 ;
        RECT 56.890 103.840 57.290 104.240 ;
        RECT 58.890 103.840 59.290 104.240 ;
        RECT 60.890 103.840 61.290 104.240 ;
        RECT 62.890 103.840 63.290 104.240 ;
        RECT 64.890 103.840 65.290 104.240 ;
        RECT 66.890 103.840 67.290 104.240 ;
        RECT 68.890 103.840 69.290 104.240 ;
        RECT 70.890 103.840 71.290 104.240 ;
        RECT 72.890 103.840 73.290 104.240 ;
        RECT 87.825 103.840 88.225 104.240 ;
        RECT 89.825 103.840 90.225 104.240 ;
        RECT 91.825 103.840 92.225 104.240 ;
        RECT 93.825 103.840 94.225 104.240 ;
        RECT 95.825 103.840 96.225 104.240 ;
        RECT 97.825 103.840 98.225 104.240 ;
        RECT 99.825 103.840 100.225 104.240 ;
        RECT 101.825 103.840 102.225 104.240 ;
        RECT 103.825 103.840 104.225 104.240 ;
        RECT 105.825 103.840 106.225 104.240 ;
        RECT 107.825 103.840 108.225 104.240 ;
        RECT 109.825 103.840 110.225 104.240 ;
        RECT 111.825 103.840 112.225 104.240 ;
        RECT 113.825 103.840 114.225 104.240 ;
        RECT 115.825 103.840 116.225 104.240 ;
        RECT 117.825 103.840 118.225 104.240 ;
        RECT 119.825 103.840 120.225 104.240 ;
        RECT 121.825 103.840 122.225 104.240 ;
        RECT 123.825 103.840 124.225 104.240 ;
        RECT 125.825 103.840 126.225 104.240 ;
        RECT 127.825 103.840 128.225 104.240 ;
        RECT 129.825 103.840 130.225 104.240 ;
        RECT 131.825 103.840 132.225 104.240 ;
        RECT 133.825 103.840 134.225 104.240 ;
        RECT 135.825 103.840 136.225 104.240 ;
        RECT 137.825 103.840 138.225 104.240 ;
        RECT 139.825 103.840 140.225 104.240 ;
        RECT 141.825 103.840 142.225 104.240 ;
        RECT 143.825 103.840 144.225 104.240 ;
        RECT 145.825 103.840 146.225 104.240 ;
        RECT 147.825 103.840 148.225 104.240 ;
        RECT 149.825 103.840 150.225 104.240 ;
        RECT 151.825 103.840 152.225 104.240 ;
        RECT 153.825 103.840 154.225 104.240 ;
        RECT 6.890 103.640 8.540 103.840 ;
        RECT 8.890 103.640 24.540 103.840 ;
        RECT 24.890 103.640 74.540 103.840 ;
        RECT 86.575 103.640 136.225 103.840 ;
        RECT 136.575 103.640 152.225 103.840 ;
        RECT 152.575 103.640 154.225 103.840 ;
        RECT 6.890 103.240 7.290 103.640 ;
        RECT 8.890 103.240 9.290 103.640 ;
        RECT 10.890 103.240 11.290 103.640 ;
        RECT 12.890 103.240 13.290 103.640 ;
        RECT 14.890 103.240 15.290 103.640 ;
        RECT 16.890 103.240 17.290 103.640 ;
        RECT 18.890 103.240 19.290 103.640 ;
        RECT 20.890 103.240 21.290 103.640 ;
        RECT 22.890 103.240 23.290 103.640 ;
        RECT 24.890 103.240 25.290 103.640 ;
        RECT 26.890 103.240 27.290 103.640 ;
        RECT 28.890 103.240 29.290 103.640 ;
        RECT 30.890 103.240 31.290 103.640 ;
        RECT 32.890 103.240 33.290 103.640 ;
        RECT 34.890 103.240 35.290 103.640 ;
        RECT 36.890 103.240 37.290 103.640 ;
        RECT 38.890 103.240 39.290 103.640 ;
        RECT 40.890 103.240 41.290 103.640 ;
        RECT 42.890 103.240 43.290 103.640 ;
        RECT 44.890 103.240 45.290 103.640 ;
        RECT 46.890 103.240 47.290 103.640 ;
        RECT 48.890 103.240 49.290 103.640 ;
        RECT 50.890 103.240 51.290 103.640 ;
        RECT 52.890 103.240 53.290 103.640 ;
        RECT 54.890 103.240 55.290 103.640 ;
        RECT 56.890 103.240 57.290 103.640 ;
        RECT 58.890 103.240 59.290 103.640 ;
        RECT 60.890 103.240 61.290 103.640 ;
        RECT 62.890 103.240 63.290 103.640 ;
        RECT 64.890 103.240 65.290 103.640 ;
        RECT 66.890 103.240 67.290 103.640 ;
        RECT 68.890 103.240 69.290 103.640 ;
        RECT 70.890 103.240 71.290 103.640 ;
        RECT 72.890 103.240 73.290 103.640 ;
        RECT 87.825 103.240 88.225 103.640 ;
        RECT 89.825 103.240 90.225 103.640 ;
        RECT 91.825 103.240 92.225 103.640 ;
        RECT 93.825 103.240 94.225 103.640 ;
        RECT 95.825 103.240 96.225 103.640 ;
        RECT 97.825 103.240 98.225 103.640 ;
        RECT 99.825 103.240 100.225 103.640 ;
        RECT 101.825 103.240 102.225 103.640 ;
        RECT 103.825 103.240 104.225 103.640 ;
        RECT 105.825 103.240 106.225 103.640 ;
        RECT 107.825 103.240 108.225 103.640 ;
        RECT 109.825 103.240 110.225 103.640 ;
        RECT 111.825 103.240 112.225 103.640 ;
        RECT 113.825 103.240 114.225 103.640 ;
        RECT 115.825 103.240 116.225 103.640 ;
        RECT 117.825 103.240 118.225 103.640 ;
        RECT 119.825 103.240 120.225 103.640 ;
        RECT 121.825 103.240 122.225 103.640 ;
        RECT 123.825 103.240 124.225 103.640 ;
        RECT 125.825 103.240 126.225 103.640 ;
        RECT 127.825 103.240 128.225 103.640 ;
        RECT 129.825 103.240 130.225 103.640 ;
        RECT 131.825 103.240 132.225 103.640 ;
        RECT 133.825 103.240 134.225 103.640 ;
        RECT 135.825 103.240 136.225 103.640 ;
        RECT 137.825 103.240 138.225 103.640 ;
        RECT 139.825 103.240 140.225 103.640 ;
        RECT 141.825 103.240 142.225 103.640 ;
        RECT 143.825 103.240 144.225 103.640 ;
        RECT 145.825 103.240 146.225 103.640 ;
        RECT 147.825 103.240 148.225 103.640 ;
        RECT 149.825 103.240 150.225 103.640 ;
        RECT 151.825 103.240 152.225 103.640 ;
        RECT 153.825 103.240 154.225 103.640 ;
        RECT 6.960 102.390 7.220 103.240 ;
        RECT 8.990 102.390 9.190 103.240 ;
        RECT 10.990 102.390 11.190 103.240 ;
        RECT 12.990 102.390 13.190 103.240 ;
        RECT 14.990 102.390 15.190 103.240 ;
        RECT 16.990 102.390 17.190 103.240 ;
        RECT 18.990 102.390 19.190 103.240 ;
        RECT 20.990 102.390 21.190 103.240 ;
        RECT 22.990 102.390 23.190 103.240 ;
        RECT 24.990 102.390 25.190 103.240 ;
        RECT 26.990 102.390 27.190 103.240 ;
        RECT 28.990 102.390 29.190 103.240 ;
        RECT 30.990 102.390 31.190 103.240 ;
        RECT 32.990 102.390 33.190 103.240 ;
        RECT 34.990 102.390 35.190 103.240 ;
        RECT 36.990 102.390 37.190 103.240 ;
        RECT 38.990 102.390 39.190 103.240 ;
        RECT 40.990 102.390 41.190 103.240 ;
        RECT 42.990 102.390 43.190 103.240 ;
        RECT 44.990 102.390 45.190 103.240 ;
        RECT 46.990 102.390 47.190 103.240 ;
        RECT 48.990 102.390 49.190 103.240 ;
        RECT 50.990 102.390 51.190 103.240 ;
        RECT 52.990 102.390 53.190 103.240 ;
        RECT 54.990 102.390 55.190 103.240 ;
        RECT 56.990 102.390 57.190 103.240 ;
        RECT 58.990 102.390 59.190 103.240 ;
        RECT 60.990 102.390 61.190 103.240 ;
        RECT 62.990 102.390 63.190 103.240 ;
        RECT 64.990 102.390 65.190 103.240 ;
        RECT 66.990 102.390 67.190 103.240 ;
        RECT 68.990 102.390 69.190 103.240 ;
        RECT 70.990 102.390 71.190 103.240 ;
        RECT 89.925 102.390 90.125 103.240 ;
        RECT 91.925 102.390 92.125 103.240 ;
        RECT 93.925 102.390 94.125 103.240 ;
        RECT 95.925 102.390 96.125 103.240 ;
        RECT 97.925 102.390 98.125 103.240 ;
        RECT 99.925 102.390 100.125 103.240 ;
        RECT 101.925 102.390 102.125 103.240 ;
        RECT 103.925 102.390 104.125 103.240 ;
        RECT 105.925 102.390 106.125 103.240 ;
        RECT 107.925 102.390 108.125 103.240 ;
        RECT 109.925 102.390 110.125 103.240 ;
        RECT 111.925 102.390 112.125 103.240 ;
        RECT 113.925 102.390 114.125 103.240 ;
        RECT 115.925 102.390 116.125 103.240 ;
        RECT 117.925 102.390 118.125 103.240 ;
        RECT 119.925 102.390 120.125 103.240 ;
        RECT 121.925 102.390 122.125 103.240 ;
        RECT 123.925 102.390 124.125 103.240 ;
        RECT 125.925 102.390 126.125 103.240 ;
        RECT 127.925 102.390 128.125 103.240 ;
        RECT 129.925 102.390 130.125 103.240 ;
        RECT 131.925 102.390 132.125 103.240 ;
        RECT 133.925 102.390 134.125 103.240 ;
        RECT 135.925 102.390 136.125 103.240 ;
        RECT 137.925 102.390 138.125 103.240 ;
        RECT 139.925 102.390 140.125 103.240 ;
        RECT 141.925 102.390 142.125 103.240 ;
        RECT 143.925 102.390 144.125 103.240 ;
        RECT 145.925 102.390 146.125 103.240 ;
        RECT 147.925 102.390 148.125 103.240 ;
        RECT 149.925 102.390 150.125 103.240 ;
        RECT 151.925 102.390 152.125 103.240 ;
        RECT 153.895 102.390 154.155 103.240 ;
        RECT 6.890 101.990 7.290 102.390 ;
        RECT 8.890 101.990 9.290 102.390 ;
        RECT 10.890 101.990 11.290 102.390 ;
        RECT 12.890 101.990 13.290 102.390 ;
        RECT 14.890 101.990 15.290 102.390 ;
        RECT 16.890 101.990 17.290 102.390 ;
        RECT 18.890 101.990 19.290 102.390 ;
        RECT 20.890 101.990 21.290 102.390 ;
        RECT 22.890 101.990 23.290 102.390 ;
        RECT 24.890 101.990 25.290 102.390 ;
        RECT 26.890 101.990 27.290 102.390 ;
        RECT 28.890 101.990 29.290 102.390 ;
        RECT 30.890 101.990 31.290 102.390 ;
        RECT 32.890 101.990 33.290 102.390 ;
        RECT 34.890 101.990 35.290 102.390 ;
        RECT 36.890 101.990 37.290 102.390 ;
        RECT 38.890 101.990 39.290 102.390 ;
        RECT 40.890 101.990 41.290 102.390 ;
        RECT 42.890 101.990 43.290 102.390 ;
        RECT 44.890 101.990 45.290 102.390 ;
        RECT 46.890 101.990 47.290 102.390 ;
        RECT 48.890 101.990 49.290 102.390 ;
        RECT 50.890 101.990 51.290 102.390 ;
        RECT 52.890 101.990 53.290 102.390 ;
        RECT 54.890 101.990 55.290 102.390 ;
        RECT 56.890 101.990 57.290 102.390 ;
        RECT 58.890 101.990 59.290 102.390 ;
        RECT 60.890 101.990 61.290 102.390 ;
        RECT 62.890 101.990 63.290 102.390 ;
        RECT 64.890 101.990 65.290 102.390 ;
        RECT 66.890 101.990 67.290 102.390 ;
        RECT 68.890 101.990 69.290 102.390 ;
        RECT 70.890 101.990 71.290 102.390 ;
        RECT 72.890 101.990 73.290 102.390 ;
        RECT 87.825 101.990 88.225 102.390 ;
        RECT 89.825 101.990 90.225 102.390 ;
        RECT 91.825 101.990 92.225 102.390 ;
        RECT 93.825 101.990 94.225 102.390 ;
        RECT 95.825 101.990 96.225 102.390 ;
        RECT 97.825 101.990 98.225 102.390 ;
        RECT 99.825 101.990 100.225 102.390 ;
        RECT 101.825 101.990 102.225 102.390 ;
        RECT 103.825 101.990 104.225 102.390 ;
        RECT 105.825 101.990 106.225 102.390 ;
        RECT 107.825 101.990 108.225 102.390 ;
        RECT 109.825 101.990 110.225 102.390 ;
        RECT 111.825 101.990 112.225 102.390 ;
        RECT 113.825 101.990 114.225 102.390 ;
        RECT 115.825 101.990 116.225 102.390 ;
        RECT 117.825 101.990 118.225 102.390 ;
        RECT 119.825 101.990 120.225 102.390 ;
        RECT 121.825 101.990 122.225 102.390 ;
        RECT 123.825 101.990 124.225 102.390 ;
        RECT 125.825 101.990 126.225 102.390 ;
        RECT 127.825 101.990 128.225 102.390 ;
        RECT 129.825 101.990 130.225 102.390 ;
        RECT 131.825 101.990 132.225 102.390 ;
        RECT 133.825 101.990 134.225 102.390 ;
        RECT 135.825 101.990 136.225 102.390 ;
        RECT 137.825 101.990 138.225 102.390 ;
        RECT 139.825 101.990 140.225 102.390 ;
        RECT 141.825 101.990 142.225 102.390 ;
        RECT 143.825 101.990 144.225 102.390 ;
        RECT 145.825 101.990 146.225 102.390 ;
        RECT 147.825 101.990 148.225 102.390 ;
        RECT 149.825 101.990 150.225 102.390 ;
        RECT 151.825 101.990 152.225 102.390 ;
        RECT 153.825 101.990 154.225 102.390 ;
        RECT 6.890 101.790 8.540 101.990 ;
        RECT 8.890 101.790 24.540 101.990 ;
        RECT 24.890 101.790 74.540 101.990 ;
        RECT 86.575 101.790 136.225 101.990 ;
        RECT 136.575 101.790 152.225 101.990 ;
        RECT 152.575 101.790 154.225 101.990 ;
        RECT 6.890 101.390 7.290 101.790 ;
        RECT 8.890 101.390 9.290 101.790 ;
        RECT 10.890 101.390 11.290 101.790 ;
        RECT 12.890 101.390 13.290 101.790 ;
        RECT 14.890 101.390 15.290 101.790 ;
        RECT 16.890 101.390 17.290 101.790 ;
        RECT 18.890 101.390 19.290 101.790 ;
        RECT 20.890 101.390 21.290 101.790 ;
        RECT 22.890 101.390 23.290 101.790 ;
        RECT 24.890 101.390 25.290 101.790 ;
        RECT 26.890 101.390 27.290 101.790 ;
        RECT 28.890 101.390 29.290 101.790 ;
        RECT 30.890 101.390 31.290 101.790 ;
        RECT 32.890 101.390 33.290 101.790 ;
        RECT 34.890 101.390 35.290 101.790 ;
        RECT 36.890 101.390 37.290 101.790 ;
        RECT 38.890 101.390 39.290 101.790 ;
        RECT 40.890 101.390 41.290 101.790 ;
        RECT 42.890 101.390 43.290 101.790 ;
        RECT 44.890 101.390 45.290 101.790 ;
        RECT 46.890 101.390 47.290 101.790 ;
        RECT 48.890 101.390 49.290 101.790 ;
        RECT 50.890 101.390 51.290 101.790 ;
        RECT 52.890 101.390 53.290 101.790 ;
        RECT 54.890 101.390 55.290 101.790 ;
        RECT 56.890 101.390 57.290 101.790 ;
        RECT 58.890 101.390 59.290 101.790 ;
        RECT 60.890 101.390 61.290 101.790 ;
        RECT 62.890 101.390 63.290 101.790 ;
        RECT 64.890 101.390 65.290 101.790 ;
        RECT 66.890 101.390 67.290 101.790 ;
        RECT 68.890 101.390 69.290 101.790 ;
        RECT 70.890 101.390 71.290 101.790 ;
        RECT 72.890 101.390 73.290 101.790 ;
        RECT 87.825 101.390 88.225 101.790 ;
        RECT 89.825 101.390 90.225 101.790 ;
        RECT 91.825 101.390 92.225 101.790 ;
        RECT 93.825 101.390 94.225 101.790 ;
        RECT 95.825 101.390 96.225 101.790 ;
        RECT 97.825 101.390 98.225 101.790 ;
        RECT 99.825 101.390 100.225 101.790 ;
        RECT 101.825 101.390 102.225 101.790 ;
        RECT 103.825 101.390 104.225 101.790 ;
        RECT 105.825 101.390 106.225 101.790 ;
        RECT 107.825 101.390 108.225 101.790 ;
        RECT 109.825 101.390 110.225 101.790 ;
        RECT 111.825 101.390 112.225 101.790 ;
        RECT 113.825 101.390 114.225 101.790 ;
        RECT 115.825 101.390 116.225 101.790 ;
        RECT 117.825 101.390 118.225 101.790 ;
        RECT 119.825 101.390 120.225 101.790 ;
        RECT 121.825 101.390 122.225 101.790 ;
        RECT 123.825 101.390 124.225 101.790 ;
        RECT 125.825 101.390 126.225 101.790 ;
        RECT 127.825 101.390 128.225 101.790 ;
        RECT 129.825 101.390 130.225 101.790 ;
        RECT 131.825 101.390 132.225 101.790 ;
        RECT 133.825 101.390 134.225 101.790 ;
        RECT 135.825 101.390 136.225 101.790 ;
        RECT 137.825 101.390 138.225 101.790 ;
        RECT 139.825 101.390 140.225 101.790 ;
        RECT 141.825 101.390 142.225 101.790 ;
        RECT 143.825 101.390 144.225 101.790 ;
        RECT 145.825 101.390 146.225 101.790 ;
        RECT 147.825 101.390 148.225 101.790 ;
        RECT 149.825 101.390 150.225 101.790 ;
        RECT 151.825 101.390 152.225 101.790 ;
        RECT 153.825 101.390 154.225 101.790 ;
        RECT 6.960 100.540 7.220 101.390 ;
        RECT 8.990 100.540 9.190 101.390 ;
        RECT 10.990 100.540 11.190 101.390 ;
        RECT 12.990 100.540 13.190 101.390 ;
        RECT 14.990 100.540 15.190 101.390 ;
        RECT 16.990 100.540 17.190 101.390 ;
        RECT 18.990 100.540 19.190 101.390 ;
        RECT 20.990 100.540 21.190 101.390 ;
        RECT 22.990 100.540 23.190 101.390 ;
        RECT 24.990 100.540 25.190 101.390 ;
        RECT 26.990 100.540 27.190 101.390 ;
        RECT 28.990 100.540 29.190 101.390 ;
        RECT 30.990 100.540 31.190 101.390 ;
        RECT 32.990 100.540 33.190 101.390 ;
        RECT 34.990 100.540 35.190 101.390 ;
        RECT 36.990 100.540 37.190 101.390 ;
        RECT 38.990 100.540 39.190 101.390 ;
        RECT 40.990 100.540 41.190 101.390 ;
        RECT 42.990 100.540 43.190 101.390 ;
        RECT 44.990 100.540 45.190 101.390 ;
        RECT 46.990 100.540 47.190 101.390 ;
        RECT 48.990 100.540 49.190 101.390 ;
        RECT 50.990 100.540 51.190 101.390 ;
        RECT 52.990 100.540 53.190 101.390 ;
        RECT 54.990 100.540 55.190 101.390 ;
        RECT 56.990 100.540 57.190 101.390 ;
        RECT 58.990 100.540 59.190 101.390 ;
        RECT 60.990 100.540 61.190 101.390 ;
        RECT 62.990 100.540 63.190 101.390 ;
        RECT 64.990 100.540 65.190 101.390 ;
        RECT 66.990 100.540 67.190 101.390 ;
        RECT 68.990 100.540 69.190 101.390 ;
        RECT 70.990 100.540 71.190 101.390 ;
        RECT 89.925 100.540 90.125 101.390 ;
        RECT 91.925 100.540 92.125 101.390 ;
        RECT 93.925 100.540 94.125 101.390 ;
        RECT 95.925 100.540 96.125 101.390 ;
        RECT 97.925 100.540 98.125 101.390 ;
        RECT 99.925 100.540 100.125 101.390 ;
        RECT 101.925 100.540 102.125 101.390 ;
        RECT 103.925 100.540 104.125 101.390 ;
        RECT 105.925 100.540 106.125 101.390 ;
        RECT 107.925 100.540 108.125 101.390 ;
        RECT 109.925 100.540 110.125 101.390 ;
        RECT 111.925 100.540 112.125 101.390 ;
        RECT 113.925 100.540 114.125 101.390 ;
        RECT 115.925 100.540 116.125 101.390 ;
        RECT 117.925 100.540 118.125 101.390 ;
        RECT 119.925 100.540 120.125 101.390 ;
        RECT 121.925 100.540 122.125 101.390 ;
        RECT 123.925 100.540 124.125 101.390 ;
        RECT 125.925 100.540 126.125 101.390 ;
        RECT 127.925 100.540 128.125 101.390 ;
        RECT 129.925 100.540 130.125 101.390 ;
        RECT 131.925 100.540 132.125 101.390 ;
        RECT 133.925 100.540 134.125 101.390 ;
        RECT 135.925 100.540 136.125 101.390 ;
        RECT 137.925 100.540 138.125 101.390 ;
        RECT 139.925 100.540 140.125 101.390 ;
        RECT 141.925 100.540 142.125 101.390 ;
        RECT 143.925 100.540 144.125 101.390 ;
        RECT 145.925 100.540 146.125 101.390 ;
        RECT 147.925 100.540 148.125 101.390 ;
        RECT 149.925 100.540 150.125 101.390 ;
        RECT 151.925 100.540 152.125 101.390 ;
        RECT 153.895 100.540 154.155 101.390 ;
        RECT 6.890 100.140 7.290 100.540 ;
        RECT 8.890 100.140 9.290 100.540 ;
        RECT 10.890 100.140 11.290 100.540 ;
        RECT 12.890 100.140 13.290 100.540 ;
        RECT 14.890 100.140 15.290 100.540 ;
        RECT 16.890 100.140 17.290 100.540 ;
        RECT 18.890 100.140 19.290 100.540 ;
        RECT 20.890 100.140 21.290 100.540 ;
        RECT 22.890 100.140 23.290 100.540 ;
        RECT 24.890 100.140 25.290 100.540 ;
        RECT 26.890 100.140 27.290 100.540 ;
        RECT 28.890 100.140 29.290 100.540 ;
        RECT 30.890 100.140 31.290 100.540 ;
        RECT 32.890 100.140 33.290 100.540 ;
        RECT 34.890 100.140 35.290 100.540 ;
        RECT 36.890 100.140 37.290 100.540 ;
        RECT 38.890 100.140 39.290 100.540 ;
        RECT 40.890 100.140 41.290 100.540 ;
        RECT 42.890 100.140 43.290 100.540 ;
        RECT 44.890 100.140 45.290 100.540 ;
        RECT 46.890 100.140 47.290 100.540 ;
        RECT 48.890 100.140 49.290 100.540 ;
        RECT 50.890 100.140 51.290 100.540 ;
        RECT 52.890 100.140 53.290 100.540 ;
        RECT 54.890 100.140 55.290 100.540 ;
        RECT 56.890 100.140 57.290 100.540 ;
        RECT 58.890 100.140 59.290 100.540 ;
        RECT 60.890 100.140 61.290 100.540 ;
        RECT 62.890 100.140 63.290 100.540 ;
        RECT 64.890 100.140 65.290 100.540 ;
        RECT 66.890 100.140 67.290 100.540 ;
        RECT 68.890 100.140 69.290 100.540 ;
        RECT 70.890 100.140 71.290 100.540 ;
        RECT 72.890 100.140 73.290 100.540 ;
        RECT 87.825 100.140 88.225 100.540 ;
        RECT 89.825 100.140 90.225 100.540 ;
        RECT 91.825 100.140 92.225 100.540 ;
        RECT 93.825 100.140 94.225 100.540 ;
        RECT 95.825 100.140 96.225 100.540 ;
        RECT 97.825 100.140 98.225 100.540 ;
        RECT 99.825 100.140 100.225 100.540 ;
        RECT 101.825 100.140 102.225 100.540 ;
        RECT 103.825 100.140 104.225 100.540 ;
        RECT 105.825 100.140 106.225 100.540 ;
        RECT 107.825 100.140 108.225 100.540 ;
        RECT 109.825 100.140 110.225 100.540 ;
        RECT 111.825 100.140 112.225 100.540 ;
        RECT 113.825 100.140 114.225 100.540 ;
        RECT 115.825 100.140 116.225 100.540 ;
        RECT 117.825 100.140 118.225 100.540 ;
        RECT 119.825 100.140 120.225 100.540 ;
        RECT 121.825 100.140 122.225 100.540 ;
        RECT 123.825 100.140 124.225 100.540 ;
        RECT 125.825 100.140 126.225 100.540 ;
        RECT 127.825 100.140 128.225 100.540 ;
        RECT 129.825 100.140 130.225 100.540 ;
        RECT 131.825 100.140 132.225 100.540 ;
        RECT 133.825 100.140 134.225 100.540 ;
        RECT 135.825 100.140 136.225 100.540 ;
        RECT 137.825 100.140 138.225 100.540 ;
        RECT 139.825 100.140 140.225 100.540 ;
        RECT 141.825 100.140 142.225 100.540 ;
        RECT 143.825 100.140 144.225 100.540 ;
        RECT 145.825 100.140 146.225 100.540 ;
        RECT 147.825 100.140 148.225 100.540 ;
        RECT 149.825 100.140 150.225 100.540 ;
        RECT 151.825 100.140 152.225 100.540 ;
        RECT 153.825 100.140 154.225 100.540 ;
        RECT 6.890 99.940 8.540 100.140 ;
        RECT 8.890 99.940 24.540 100.140 ;
        RECT 24.890 99.940 74.540 100.140 ;
        RECT 86.575 99.940 136.225 100.140 ;
        RECT 136.575 99.940 152.225 100.140 ;
        RECT 152.575 99.940 154.225 100.140 ;
        RECT 6.890 99.540 7.290 99.940 ;
        RECT 8.890 99.540 9.290 99.940 ;
        RECT 10.890 99.540 11.290 99.940 ;
        RECT 12.890 99.540 13.290 99.940 ;
        RECT 14.890 99.540 15.290 99.940 ;
        RECT 16.890 99.540 17.290 99.940 ;
        RECT 18.890 99.540 19.290 99.940 ;
        RECT 20.890 99.540 21.290 99.940 ;
        RECT 22.890 99.540 23.290 99.940 ;
        RECT 24.890 99.540 25.290 99.940 ;
        RECT 26.890 99.540 27.290 99.940 ;
        RECT 28.890 99.540 29.290 99.940 ;
        RECT 30.890 99.540 31.290 99.940 ;
        RECT 32.890 99.540 33.290 99.940 ;
        RECT 34.890 99.540 35.290 99.940 ;
        RECT 36.890 99.540 37.290 99.940 ;
        RECT 38.890 99.540 39.290 99.940 ;
        RECT 40.890 99.540 41.290 99.940 ;
        RECT 42.890 99.540 43.290 99.940 ;
        RECT 44.890 99.540 45.290 99.940 ;
        RECT 46.890 99.540 47.290 99.940 ;
        RECT 48.890 99.540 49.290 99.940 ;
        RECT 50.890 99.540 51.290 99.940 ;
        RECT 52.890 99.540 53.290 99.940 ;
        RECT 54.890 99.540 55.290 99.940 ;
        RECT 56.890 99.540 57.290 99.940 ;
        RECT 58.890 99.540 59.290 99.940 ;
        RECT 60.890 99.540 61.290 99.940 ;
        RECT 62.890 99.540 63.290 99.940 ;
        RECT 64.890 99.540 65.290 99.940 ;
        RECT 66.890 99.540 67.290 99.940 ;
        RECT 68.890 99.540 69.290 99.940 ;
        RECT 70.890 99.540 71.290 99.940 ;
        RECT 72.890 99.540 73.290 99.940 ;
        RECT 87.825 99.540 88.225 99.940 ;
        RECT 89.825 99.540 90.225 99.940 ;
        RECT 91.825 99.540 92.225 99.940 ;
        RECT 93.825 99.540 94.225 99.940 ;
        RECT 95.825 99.540 96.225 99.940 ;
        RECT 97.825 99.540 98.225 99.940 ;
        RECT 99.825 99.540 100.225 99.940 ;
        RECT 101.825 99.540 102.225 99.940 ;
        RECT 103.825 99.540 104.225 99.940 ;
        RECT 105.825 99.540 106.225 99.940 ;
        RECT 107.825 99.540 108.225 99.940 ;
        RECT 109.825 99.540 110.225 99.940 ;
        RECT 111.825 99.540 112.225 99.940 ;
        RECT 113.825 99.540 114.225 99.940 ;
        RECT 115.825 99.540 116.225 99.940 ;
        RECT 117.825 99.540 118.225 99.940 ;
        RECT 119.825 99.540 120.225 99.940 ;
        RECT 121.825 99.540 122.225 99.940 ;
        RECT 123.825 99.540 124.225 99.940 ;
        RECT 125.825 99.540 126.225 99.940 ;
        RECT 127.825 99.540 128.225 99.940 ;
        RECT 129.825 99.540 130.225 99.940 ;
        RECT 131.825 99.540 132.225 99.940 ;
        RECT 133.825 99.540 134.225 99.940 ;
        RECT 135.825 99.540 136.225 99.940 ;
        RECT 137.825 99.540 138.225 99.940 ;
        RECT 139.825 99.540 140.225 99.940 ;
        RECT 141.825 99.540 142.225 99.940 ;
        RECT 143.825 99.540 144.225 99.940 ;
        RECT 145.825 99.540 146.225 99.940 ;
        RECT 147.825 99.540 148.225 99.940 ;
        RECT 149.825 99.540 150.225 99.940 ;
        RECT 151.825 99.540 152.225 99.940 ;
        RECT 153.825 99.540 154.225 99.940 ;
        RECT 6.960 98.690 7.220 99.540 ;
        RECT 8.990 98.690 9.190 99.540 ;
        RECT 10.990 98.690 11.190 99.540 ;
        RECT 12.990 98.690 13.190 99.540 ;
        RECT 14.990 98.690 15.190 99.540 ;
        RECT 16.990 98.690 17.190 99.540 ;
        RECT 18.990 98.690 19.190 99.540 ;
        RECT 20.990 98.690 21.190 99.540 ;
        RECT 22.990 98.690 23.190 99.540 ;
        RECT 24.990 98.690 25.190 99.540 ;
        RECT 26.990 98.690 27.190 99.540 ;
        RECT 28.990 98.690 29.190 99.540 ;
        RECT 30.990 98.690 31.190 99.540 ;
        RECT 32.990 98.690 33.190 99.540 ;
        RECT 34.990 98.690 35.190 99.540 ;
        RECT 36.990 98.690 37.190 99.540 ;
        RECT 38.990 98.690 39.190 99.540 ;
        RECT 40.990 98.690 41.190 99.540 ;
        RECT 42.990 98.690 43.190 99.540 ;
        RECT 44.990 98.690 45.190 99.540 ;
        RECT 46.990 98.690 47.190 99.540 ;
        RECT 48.990 98.690 49.190 99.540 ;
        RECT 50.990 98.690 51.190 99.540 ;
        RECT 52.990 98.690 53.190 99.540 ;
        RECT 54.990 98.690 55.190 99.540 ;
        RECT 56.990 98.690 57.190 99.540 ;
        RECT 58.990 98.690 59.190 99.540 ;
        RECT 60.990 98.690 61.190 99.540 ;
        RECT 62.990 98.690 63.190 99.540 ;
        RECT 64.990 98.690 65.190 99.540 ;
        RECT 66.990 98.690 67.190 99.540 ;
        RECT 68.990 98.690 69.190 99.540 ;
        RECT 70.990 98.690 71.190 99.540 ;
        RECT 89.925 98.690 90.125 99.540 ;
        RECT 91.925 98.690 92.125 99.540 ;
        RECT 93.925 98.690 94.125 99.540 ;
        RECT 95.925 98.690 96.125 99.540 ;
        RECT 97.925 98.690 98.125 99.540 ;
        RECT 99.925 98.690 100.125 99.540 ;
        RECT 101.925 98.690 102.125 99.540 ;
        RECT 103.925 98.690 104.125 99.540 ;
        RECT 105.925 98.690 106.125 99.540 ;
        RECT 107.925 98.690 108.125 99.540 ;
        RECT 109.925 98.690 110.125 99.540 ;
        RECT 111.925 98.690 112.125 99.540 ;
        RECT 113.925 98.690 114.125 99.540 ;
        RECT 115.925 98.690 116.125 99.540 ;
        RECT 117.925 98.690 118.125 99.540 ;
        RECT 119.925 98.690 120.125 99.540 ;
        RECT 121.925 98.690 122.125 99.540 ;
        RECT 123.925 98.690 124.125 99.540 ;
        RECT 125.925 98.690 126.125 99.540 ;
        RECT 127.925 98.690 128.125 99.540 ;
        RECT 129.925 98.690 130.125 99.540 ;
        RECT 131.925 98.690 132.125 99.540 ;
        RECT 133.925 98.690 134.125 99.540 ;
        RECT 135.925 98.690 136.125 99.540 ;
        RECT 137.925 98.690 138.125 99.540 ;
        RECT 139.925 98.690 140.125 99.540 ;
        RECT 141.925 98.690 142.125 99.540 ;
        RECT 143.925 98.690 144.125 99.540 ;
        RECT 145.925 98.690 146.125 99.540 ;
        RECT 147.925 98.690 148.125 99.540 ;
        RECT 149.925 98.690 150.125 99.540 ;
        RECT 151.925 98.690 152.125 99.540 ;
        RECT 153.895 98.690 154.155 99.540 ;
        RECT 6.890 98.290 7.290 98.690 ;
        RECT 8.890 98.290 9.290 98.690 ;
        RECT 10.890 98.290 11.290 98.690 ;
        RECT 12.890 98.290 13.290 98.690 ;
        RECT 14.890 98.290 15.290 98.690 ;
        RECT 16.890 98.290 17.290 98.690 ;
        RECT 18.890 98.290 19.290 98.690 ;
        RECT 20.890 98.290 21.290 98.690 ;
        RECT 22.890 98.290 23.290 98.690 ;
        RECT 24.890 98.290 25.290 98.690 ;
        RECT 26.890 98.290 27.290 98.690 ;
        RECT 28.890 98.290 29.290 98.690 ;
        RECT 30.890 98.290 31.290 98.690 ;
        RECT 32.890 98.290 33.290 98.690 ;
        RECT 34.890 98.290 35.290 98.690 ;
        RECT 36.890 98.290 37.290 98.690 ;
        RECT 38.890 98.290 39.290 98.690 ;
        RECT 40.890 98.290 41.290 98.690 ;
        RECT 42.890 98.290 43.290 98.690 ;
        RECT 44.890 98.290 45.290 98.690 ;
        RECT 46.890 98.290 47.290 98.690 ;
        RECT 48.890 98.290 49.290 98.690 ;
        RECT 50.890 98.290 51.290 98.690 ;
        RECT 52.890 98.290 53.290 98.690 ;
        RECT 54.890 98.290 55.290 98.690 ;
        RECT 56.890 98.290 57.290 98.690 ;
        RECT 58.890 98.290 59.290 98.690 ;
        RECT 60.890 98.290 61.290 98.690 ;
        RECT 62.890 98.290 63.290 98.690 ;
        RECT 64.890 98.290 65.290 98.690 ;
        RECT 66.890 98.290 67.290 98.690 ;
        RECT 68.890 98.290 69.290 98.690 ;
        RECT 70.890 98.290 71.290 98.690 ;
        RECT 72.890 98.290 73.290 98.690 ;
        RECT 87.825 98.290 88.225 98.690 ;
        RECT 89.825 98.290 90.225 98.690 ;
        RECT 91.825 98.290 92.225 98.690 ;
        RECT 93.825 98.290 94.225 98.690 ;
        RECT 95.825 98.290 96.225 98.690 ;
        RECT 97.825 98.290 98.225 98.690 ;
        RECT 99.825 98.290 100.225 98.690 ;
        RECT 101.825 98.290 102.225 98.690 ;
        RECT 103.825 98.290 104.225 98.690 ;
        RECT 105.825 98.290 106.225 98.690 ;
        RECT 107.825 98.290 108.225 98.690 ;
        RECT 109.825 98.290 110.225 98.690 ;
        RECT 111.825 98.290 112.225 98.690 ;
        RECT 113.825 98.290 114.225 98.690 ;
        RECT 115.825 98.290 116.225 98.690 ;
        RECT 117.825 98.290 118.225 98.690 ;
        RECT 119.825 98.290 120.225 98.690 ;
        RECT 121.825 98.290 122.225 98.690 ;
        RECT 123.825 98.290 124.225 98.690 ;
        RECT 125.825 98.290 126.225 98.690 ;
        RECT 127.825 98.290 128.225 98.690 ;
        RECT 129.825 98.290 130.225 98.690 ;
        RECT 131.825 98.290 132.225 98.690 ;
        RECT 133.825 98.290 134.225 98.690 ;
        RECT 135.825 98.290 136.225 98.690 ;
        RECT 137.825 98.290 138.225 98.690 ;
        RECT 139.825 98.290 140.225 98.690 ;
        RECT 141.825 98.290 142.225 98.690 ;
        RECT 143.825 98.290 144.225 98.690 ;
        RECT 145.825 98.290 146.225 98.690 ;
        RECT 147.825 98.290 148.225 98.690 ;
        RECT 149.825 98.290 150.225 98.690 ;
        RECT 151.825 98.290 152.225 98.690 ;
        RECT 153.825 98.290 154.225 98.690 ;
        RECT 6.890 98.090 8.540 98.290 ;
        RECT 8.890 98.090 24.540 98.290 ;
        RECT 24.890 98.090 74.540 98.290 ;
        RECT 86.575 98.090 136.225 98.290 ;
        RECT 136.575 98.090 152.225 98.290 ;
        RECT 152.575 98.090 154.225 98.290 ;
        RECT 6.890 97.690 7.290 98.090 ;
        RECT 8.890 97.690 9.290 98.090 ;
        RECT 10.890 97.690 11.290 98.090 ;
        RECT 12.890 97.690 13.290 98.090 ;
        RECT 14.890 97.690 15.290 98.090 ;
        RECT 16.890 97.690 17.290 98.090 ;
        RECT 18.890 97.690 19.290 98.090 ;
        RECT 20.890 97.690 21.290 98.090 ;
        RECT 22.890 97.690 23.290 98.090 ;
        RECT 24.890 97.690 25.290 98.090 ;
        RECT 26.890 97.690 27.290 98.090 ;
        RECT 28.890 97.690 29.290 98.090 ;
        RECT 30.890 97.690 31.290 98.090 ;
        RECT 32.890 97.690 33.290 98.090 ;
        RECT 34.890 97.690 35.290 98.090 ;
        RECT 36.890 97.690 37.290 98.090 ;
        RECT 38.890 97.690 39.290 98.090 ;
        RECT 40.890 97.690 41.290 98.090 ;
        RECT 42.890 97.690 43.290 98.090 ;
        RECT 44.890 97.690 45.290 98.090 ;
        RECT 46.890 97.690 47.290 98.090 ;
        RECT 48.890 97.690 49.290 98.090 ;
        RECT 50.890 97.690 51.290 98.090 ;
        RECT 52.890 97.690 53.290 98.090 ;
        RECT 54.890 97.690 55.290 98.090 ;
        RECT 56.890 97.690 57.290 98.090 ;
        RECT 58.890 97.690 59.290 98.090 ;
        RECT 60.890 97.690 61.290 98.090 ;
        RECT 62.890 97.690 63.290 98.090 ;
        RECT 64.890 97.690 65.290 98.090 ;
        RECT 66.890 97.690 67.290 98.090 ;
        RECT 68.890 97.690 69.290 98.090 ;
        RECT 70.890 97.690 71.290 98.090 ;
        RECT 72.890 97.690 73.290 98.090 ;
        RECT 87.825 97.690 88.225 98.090 ;
        RECT 89.825 97.690 90.225 98.090 ;
        RECT 91.825 97.690 92.225 98.090 ;
        RECT 93.825 97.690 94.225 98.090 ;
        RECT 95.825 97.690 96.225 98.090 ;
        RECT 97.825 97.690 98.225 98.090 ;
        RECT 99.825 97.690 100.225 98.090 ;
        RECT 101.825 97.690 102.225 98.090 ;
        RECT 103.825 97.690 104.225 98.090 ;
        RECT 105.825 97.690 106.225 98.090 ;
        RECT 107.825 97.690 108.225 98.090 ;
        RECT 109.825 97.690 110.225 98.090 ;
        RECT 111.825 97.690 112.225 98.090 ;
        RECT 113.825 97.690 114.225 98.090 ;
        RECT 115.825 97.690 116.225 98.090 ;
        RECT 117.825 97.690 118.225 98.090 ;
        RECT 119.825 97.690 120.225 98.090 ;
        RECT 121.825 97.690 122.225 98.090 ;
        RECT 123.825 97.690 124.225 98.090 ;
        RECT 125.825 97.690 126.225 98.090 ;
        RECT 127.825 97.690 128.225 98.090 ;
        RECT 129.825 97.690 130.225 98.090 ;
        RECT 131.825 97.690 132.225 98.090 ;
        RECT 133.825 97.690 134.225 98.090 ;
        RECT 135.825 97.690 136.225 98.090 ;
        RECT 137.825 97.690 138.225 98.090 ;
        RECT 139.825 97.690 140.225 98.090 ;
        RECT 141.825 97.690 142.225 98.090 ;
        RECT 143.825 97.690 144.225 98.090 ;
        RECT 145.825 97.690 146.225 98.090 ;
        RECT 147.825 97.690 148.225 98.090 ;
        RECT 149.825 97.690 150.225 98.090 ;
        RECT 151.825 97.690 152.225 98.090 ;
        RECT 153.825 97.690 154.225 98.090 ;
        RECT 6.960 96.840 7.220 97.690 ;
        RECT 8.990 96.840 9.190 97.690 ;
        RECT 10.990 96.840 11.190 97.690 ;
        RECT 12.990 96.840 13.190 97.690 ;
        RECT 14.990 96.840 15.190 97.690 ;
        RECT 16.990 96.840 17.190 97.690 ;
        RECT 18.990 96.840 19.190 97.690 ;
        RECT 20.990 96.840 21.190 97.690 ;
        RECT 22.990 96.840 23.190 97.690 ;
        RECT 24.990 96.840 25.190 97.690 ;
        RECT 26.990 96.840 27.190 97.690 ;
        RECT 28.990 96.840 29.190 97.690 ;
        RECT 30.990 96.840 31.190 97.690 ;
        RECT 32.990 96.840 33.190 97.690 ;
        RECT 34.990 96.840 35.190 97.690 ;
        RECT 36.990 96.840 37.190 97.690 ;
        RECT 38.990 96.840 39.190 97.690 ;
        RECT 40.990 96.840 41.190 97.690 ;
        RECT 42.990 96.840 43.190 97.690 ;
        RECT 44.990 96.840 45.190 97.690 ;
        RECT 46.990 96.840 47.190 97.690 ;
        RECT 48.990 96.840 49.190 97.690 ;
        RECT 50.990 96.840 51.190 97.690 ;
        RECT 52.990 96.840 53.190 97.690 ;
        RECT 54.990 96.840 55.190 97.690 ;
        RECT 56.990 96.840 57.190 97.690 ;
        RECT 58.990 96.840 59.190 97.690 ;
        RECT 60.990 96.840 61.190 97.690 ;
        RECT 62.990 96.840 63.190 97.690 ;
        RECT 64.990 96.840 65.190 97.690 ;
        RECT 66.990 96.840 67.190 97.690 ;
        RECT 68.990 96.840 69.190 97.690 ;
        RECT 70.990 96.840 71.190 97.690 ;
        RECT 89.925 96.840 90.125 97.690 ;
        RECT 91.925 96.840 92.125 97.690 ;
        RECT 93.925 96.840 94.125 97.690 ;
        RECT 95.925 96.840 96.125 97.690 ;
        RECT 97.925 96.840 98.125 97.690 ;
        RECT 99.925 96.840 100.125 97.690 ;
        RECT 101.925 96.840 102.125 97.690 ;
        RECT 103.925 96.840 104.125 97.690 ;
        RECT 105.925 96.840 106.125 97.690 ;
        RECT 107.925 96.840 108.125 97.690 ;
        RECT 109.925 96.840 110.125 97.690 ;
        RECT 111.925 96.840 112.125 97.690 ;
        RECT 113.925 96.840 114.125 97.690 ;
        RECT 115.925 96.840 116.125 97.690 ;
        RECT 117.925 96.840 118.125 97.690 ;
        RECT 119.925 96.840 120.125 97.690 ;
        RECT 121.925 96.840 122.125 97.690 ;
        RECT 123.925 96.840 124.125 97.690 ;
        RECT 125.925 96.840 126.125 97.690 ;
        RECT 127.925 96.840 128.125 97.690 ;
        RECT 129.925 96.840 130.125 97.690 ;
        RECT 131.925 96.840 132.125 97.690 ;
        RECT 133.925 96.840 134.125 97.690 ;
        RECT 135.925 96.840 136.125 97.690 ;
        RECT 137.925 96.840 138.125 97.690 ;
        RECT 139.925 96.840 140.125 97.690 ;
        RECT 141.925 96.840 142.125 97.690 ;
        RECT 143.925 96.840 144.125 97.690 ;
        RECT 145.925 96.840 146.125 97.690 ;
        RECT 147.925 96.840 148.125 97.690 ;
        RECT 149.925 96.840 150.125 97.690 ;
        RECT 151.925 96.840 152.125 97.690 ;
        RECT 153.895 96.840 154.155 97.690 ;
        RECT 6.890 96.440 7.290 96.840 ;
        RECT 8.890 96.440 9.290 96.840 ;
        RECT 10.890 96.440 11.290 96.840 ;
        RECT 12.890 96.440 13.290 96.840 ;
        RECT 14.890 96.440 15.290 96.840 ;
        RECT 16.890 96.440 17.290 96.840 ;
        RECT 18.890 96.440 19.290 96.840 ;
        RECT 20.890 96.440 21.290 96.840 ;
        RECT 22.890 96.440 23.290 96.840 ;
        RECT 24.890 96.440 25.290 96.840 ;
        RECT 26.890 96.440 27.290 96.840 ;
        RECT 28.890 96.440 29.290 96.840 ;
        RECT 30.890 96.440 31.290 96.840 ;
        RECT 32.890 96.440 33.290 96.840 ;
        RECT 34.890 96.440 35.290 96.840 ;
        RECT 36.890 96.440 37.290 96.840 ;
        RECT 38.890 96.440 39.290 96.840 ;
        RECT 40.890 96.440 41.290 96.840 ;
        RECT 42.890 96.440 43.290 96.840 ;
        RECT 44.890 96.440 45.290 96.840 ;
        RECT 46.890 96.440 47.290 96.840 ;
        RECT 48.890 96.440 49.290 96.840 ;
        RECT 50.890 96.440 51.290 96.840 ;
        RECT 52.890 96.440 53.290 96.840 ;
        RECT 54.890 96.440 55.290 96.840 ;
        RECT 56.890 96.440 57.290 96.840 ;
        RECT 58.890 96.440 59.290 96.840 ;
        RECT 60.890 96.440 61.290 96.840 ;
        RECT 62.890 96.440 63.290 96.840 ;
        RECT 64.890 96.440 65.290 96.840 ;
        RECT 66.890 96.440 67.290 96.840 ;
        RECT 68.890 96.440 69.290 96.840 ;
        RECT 70.890 96.440 71.290 96.840 ;
        RECT 72.890 96.440 73.290 96.840 ;
        RECT 87.825 96.440 88.225 96.840 ;
        RECT 89.825 96.440 90.225 96.840 ;
        RECT 91.825 96.440 92.225 96.840 ;
        RECT 93.825 96.440 94.225 96.840 ;
        RECT 95.825 96.440 96.225 96.840 ;
        RECT 97.825 96.440 98.225 96.840 ;
        RECT 99.825 96.440 100.225 96.840 ;
        RECT 101.825 96.440 102.225 96.840 ;
        RECT 103.825 96.440 104.225 96.840 ;
        RECT 105.825 96.440 106.225 96.840 ;
        RECT 107.825 96.440 108.225 96.840 ;
        RECT 109.825 96.440 110.225 96.840 ;
        RECT 111.825 96.440 112.225 96.840 ;
        RECT 113.825 96.440 114.225 96.840 ;
        RECT 115.825 96.440 116.225 96.840 ;
        RECT 117.825 96.440 118.225 96.840 ;
        RECT 119.825 96.440 120.225 96.840 ;
        RECT 121.825 96.440 122.225 96.840 ;
        RECT 123.825 96.440 124.225 96.840 ;
        RECT 125.825 96.440 126.225 96.840 ;
        RECT 127.825 96.440 128.225 96.840 ;
        RECT 129.825 96.440 130.225 96.840 ;
        RECT 131.825 96.440 132.225 96.840 ;
        RECT 133.825 96.440 134.225 96.840 ;
        RECT 135.825 96.440 136.225 96.840 ;
        RECT 137.825 96.440 138.225 96.840 ;
        RECT 139.825 96.440 140.225 96.840 ;
        RECT 141.825 96.440 142.225 96.840 ;
        RECT 143.825 96.440 144.225 96.840 ;
        RECT 145.825 96.440 146.225 96.840 ;
        RECT 147.825 96.440 148.225 96.840 ;
        RECT 149.825 96.440 150.225 96.840 ;
        RECT 151.825 96.440 152.225 96.840 ;
        RECT 153.825 96.440 154.225 96.840 ;
        RECT 6.890 96.240 8.540 96.440 ;
        RECT 8.890 96.240 24.540 96.440 ;
        RECT 24.890 96.240 74.540 96.440 ;
        RECT 86.575 96.240 136.225 96.440 ;
        RECT 136.575 96.240 152.225 96.440 ;
        RECT 152.575 96.240 154.225 96.440 ;
        RECT 6.890 95.840 7.290 96.240 ;
        RECT 8.890 95.840 9.290 96.240 ;
        RECT 10.890 95.840 11.290 96.240 ;
        RECT 12.890 95.840 13.290 96.240 ;
        RECT 14.890 95.840 15.290 96.240 ;
        RECT 16.890 95.840 17.290 96.240 ;
        RECT 18.890 95.840 19.290 96.240 ;
        RECT 20.890 95.840 21.290 96.240 ;
        RECT 22.890 95.840 23.290 96.240 ;
        RECT 24.890 95.840 25.290 96.240 ;
        RECT 26.890 95.840 27.290 96.240 ;
        RECT 28.890 95.840 29.290 96.240 ;
        RECT 30.890 95.840 31.290 96.240 ;
        RECT 32.890 95.840 33.290 96.240 ;
        RECT 34.890 95.840 35.290 96.240 ;
        RECT 36.890 95.840 37.290 96.240 ;
        RECT 38.890 95.840 39.290 96.240 ;
        RECT 40.890 95.840 41.290 96.240 ;
        RECT 42.890 95.840 43.290 96.240 ;
        RECT 44.890 95.840 45.290 96.240 ;
        RECT 46.890 95.840 47.290 96.240 ;
        RECT 48.890 95.840 49.290 96.240 ;
        RECT 50.890 95.840 51.290 96.240 ;
        RECT 52.890 95.840 53.290 96.240 ;
        RECT 54.890 95.840 55.290 96.240 ;
        RECT 56.890 95.840 57.290 96.240 ;
        RECT 58.890 95.840 59.290 96.240 ;
        RECT 60.890 95.840 61.290 96.240 ;
        RECT 62.890 95.840 63.290 96.240 ;
        RECT 64.890 95.840 65.290 96.240 ;
        RECT 66.890 95.840 67.290 96.240 ;
        RECT 68.890 95.840 69.290 96.240 ;
        RECT 70.890 95.840 71.290 96.240 ;
        RECT 72.890 95.840 73.290 96.240 ;
        RECT 87.825 95.840 88.225 96.240 ;
        RECT 89.825 95.840 90.225 96.240 ;
        RECT 91.825 95.840 92.225 96.240 ;
        RECT 93.825 95.840 94.225 96.240 ;
        RECT 95.825 95.840 96.225 96.240 ;
        RECT 97.825 95.840 98.225 96.240 ;
        RECT 99.825 95.840 100.225 96.240 ;
        RECT 101.825 95.840 102.225 96.240 ;
        RECT 103.825 95.840 104.225 96.240 ;
        RECT 105.825 95.840 106.225 96.240 ;
        RECT 107.825 95.840 108.225 96.240 ;
        RECT 109.825 95.840 110.225 96.240 ;
        RECT 111.825 95.840 112.225 96.240 ;
        RECT 113.825 95.840 114.225 96.240 ;
        RECT 115.825 95.840 116.225 96.240 ;
        RECT 117.825 95.840 118.225 96.240 ;
        RECT 119.825 95.840 120.225 96.240 ;
        RECT 121.825 95.840 122.225 96.240 ;
        RECT 123.825 95.840 124.225 96.240 ;
        RECT 125.825 95.840 126.225 96.240 ;
        RECT 127.825 95.840 128.225 96.240 ;
        RECT 129.825 95.840 130.225 96.240 ;
        RECT 131.825 95.840 132.225 96.240 ;
        RECT 133.825 95.840 134.225 96.240 ;
        RECT 135.825 95.840 136.225 96.240 ;
        RECT 137.825 95.840 138.225 96.240 ;
        RECT 139.825 95.840 140.225 96.240 ;
        RECT 141.825 95.840 142.225 96.240 ;
        RECT 143.825 95.840 144.225 96.240 ;
        RECT 145.825 95.840 146.225 96.240 ;
        RECT 147.825 95.840 148.225 96.240 ;
        RECT 149.825 95.840 150.225 96.240 ;
        RECT 151.825 95.840 152.225 96.240 ;
        RECT 153.825 95.840 154.225 96.240 ;
        RECT 6.960 94.990 7.220 95.840 ;
        RECT 8.990 94.990 9.190 95.840 ;
        RECT 10.990 94.990 11.190 95.840 ;
        RECT 12.990 94.990 13.190 95.840 ;
        RECT 14.990 94.990 15.190 95.840 ;
        RECT 16.990 94.990 17.190 95.840 ;
        RECT 18.990 94.990 19.190 95.840 ;
        RECT 20.990 94.990 21.190 95.840 ;
        RECT 22.990 94.990 23.190 95.840 ;
        RECT 24.990 94.990 25.190 95.840 ;
        RECT 26.990 94.990 27.190 95.840 ;
        RECT 28.990 94.990 29.190 95.840 ;
        RECT 30.990 94.990 31.190 95.840 ;
        RECT 32.990 94.990 33.190 95.840 ;
        RECT 34.990 94.990 35.190 95.840 ;
        RECT 36.990 94.990 37.190 95.840 ;
        RECT 38.990 94.990 39.190 95.840 ;
        RECT 40.990 94.990 41.190 95.840 ;
        RECT 42.990 94.990 43.190 95.840 ;
        RECT 44.990 94.990 45.190 95.840 ;
        RECT 46.990 94.990 47.190 95.840 ;
        RECT 48.990 94.990 49.190 95.840 ;
        RECT 50.990 94.990 51.190 95.840 ;
        RECT 52.990 94.990 53.190 95.840 ;
        RECT 54.990 94.990 55.190 95.840 ;
        RECT 56.990 94.990 57.190 95.840 ;
        RECT 58.990 94.990 59.190 95.840 ;
        RECT 60.990 94.990 61.190 95.840 ;
        RECT 62.990 94.990 63.190 95.840 ;
        RECT 64.990 94.990 65.190 95.840 ;
        RECT 66.990 94.990 67.190 95.840 ;
        RECT 68.990 94.990 69.190 95.840 ;
        RECT 70.990 94.990 71.190 95.840 ;
        RECT 89.925 94.990 90.125 95.840 ;
        RECT 91.925 94.990 92.125 95.840 ;
        RECT 93.925 94.990 94.125 95.840 ;
        RECT 95.925 94.990 96.125 95.840 ;
        RECT 97.925 94.990 98.125 95.840 ;
        RECT 99.925 94.990 100.125 95.840 ;
        RECT 101.925 94.990 102.125 95.840 ;
        RECT 103.925 94.990 104.125 95.840 ;
        RECT 105.925 94.990 106.125 95.840 ;
        RECT 107.925 94.990 108.125 95.840 ;
        RECT 109.925 94.990 110.125 95.840 ;
        RECT 111.925 94.990 112.125 95.840 ;
        RECT 113.925 94.990 114.125 95.840 ;
        RECT 115.925 94.990 116.125 95.840 ;
        RECT 117.925 94.990 118.125 95.840 ;
        RECT 119.925 94.990 120.125 95.840 ;
        RECT 121.925 94.990 122.125 95.840 ;
        RECT 123.925 94.990 124.125 95.840 ;
        RECT 125.925 94.990 126.125 95.840 ;
        RECT 127.925 94.990 128.125 95.840 ;
        RECT 129.925 94.990 130.125 95.840 ;
        RECT 131.925 94.990 132.125 95.840 ;
        RECT 133.925 94.990 134.125 95.840 ;
        RECT 135.925 94.990 136.125 95.840 ;
        RECT 137.925 94.990 138.125 95.840 ;
        RECT 139.925 94.990 140.125 95.840 ;
        RECT 141.925 94.990 142.125 95.840 ;
        RECT 143.925 94.990 144.125 95.840 ;
        RECT 145.925 94.990 146.125 95.840 ;
        RECT 147.925 94.990 148.125 95.840 ;
        RECT 149.925 94.990 150.125 95.840 ;
        RECT 151.925 94.990 152.125 95.840 ;
        RECT 153.895 94.990 154.155 95.840 ;
        RECT 6.890 94.590 7.290 94.990 ;
        RECT 8.890 94.590 9.290 94.990 ;
        RECT 10.890 94.590 11.290 94.990 ;
        RECT 12.890 94.590 13.290 94.990 ;
        RECT 14.890 94.590 15.290 94.990 ;
        RECT 16.890 94.590 17.290 94.990 ;
        RECT 18.890 94.590 19.290 94.990 ;
        RECT 20.890 94.590 21.290 94.990 ;
        RECT 22.890 94.590 23.290 94.990 ;
        RECT 24.890 94.590 25.290 94.990 ;
        RECT 26.890 94.590 27.290 94.990 ;
        RECT 28.890 94.590 29.290 94.990 ;
        RECT 30.890 94.590 31.290 94.990 ;
        RECT 32.890 94.590 33.290 94.990 ;
        RECT 34.890 94.590 35.290 94.990 ;
        RECT 36.890 94.590 37.290 94.990 ;
        RECT 38.890 94.590 39.290 94.990 ;
        RECT 40.890 94.590 41.290 94.990 ;
        RECT 42.890 94.590 43.290 94.990 ;
        RECT 44.890 94.590 45.290 94.990 ;
        RECT 46.890 94.590 47.290 94.990 ;
        RECT 48.890 94.590 49.290 94.990 ;
        RECT 50.890 94.590 51.290 94.990 ;
        RECT 52.890 94.590 53.290 94.990 ;
        RECT 54.890 94.590 55.290 94.990 ;
        RECT 56.890 94.590 57.290 94.990 ;
        RECT 58.890 94.590 59.290 94.990 ;
        RECT 60.890 94.590 61.290 94.990 ;
        RECT 62.890 94.590 63.290 94.990 ;
        RECT 64.890 94.590 65.290 94.990 ;
        RECT 66.890 94.590 67.290 94.990 ;
        RECT 68.890 94.590 69.290 94.990 ;
        RECT 70.890 94.590 71.290 94.990 ;
        RECT 72.890 94.590 73.290 94.990 ;
        RECT 87.825 94.590 88.225 94.990 ;
        RECT 89.825 94.590 90.225 94.990 ;
        RECT 91.825 94.590 92.225 94.990 ;
        RECT 93.825 94.590 94.225 94.990 ;
        RECT 95.825 94.590 96.225 94.990 ;
        RECT 97.825 94.590 98.225 94.990 ;
        RECT 99.825 94.590 100.225 94.990 ;
        RECT 101.825 94.590 102.225 94.990 ;
        RECT 103.825 94.590 104.225 94.990 ;
        RECT 105.825 94.590 106.225 94.990 ;
        RECT 107.825 94.590 108.225 94.990 ;
        RECT 109.825 94.590 110.225 94.990 ;
        RECT 111.825 94.590 112.225 94.990 ;
        RECT 113.825 94.590 114.225 94.990 ;
        RECT 115.825 94.590 116.225 94.990 ;
        RECT 117.825 94.590 118.225 94.990 ;
        RECT 119.825 94.590 120.225 94.990 ;
        RECT 121.825 94.590 122.225 94.990 ;
        RECT 123.825 94.590 124.225 94.990 ;
        RECT 125.825 94.590 126.225 94.990 ;
        RECT 127.825 94.590 128.225 94.990 ;
        RECT 129.825 94.590 130.225 94.990 ;
        RECT 131.825 94.590 132.225 94.990 ;
        RECT 133.825 94.590 134.225 94.990 ;
        RECT 135.825 94.590 136.225 94.990 ;
        RECT 137.825 94.590 138.225 94.990 ;
        RECT 139.825 94.590 140.225 94.990 ;
        RECT 141.825 94.590 142.225 94.990 ;
        RECT 143.825 94.590 144.225 94.990 ;
        RECT 145.825 94.590 146.225 94.990 ;
        RECT 147.825 94.590 148.225 94.990 ;
        RECT 149.825 94.590 150.225 94.990 ;
        RECT 151.825 94.590 152.225 94.990 ;
        RECT 153.825 94.590 154.225 94.990 ;
        RECT 6.890 94.390 8.540 94.590 ;
        RECT 8.890 94.390 24.540 94.590 ;
        RECT 24.890 94.390 74.540 94.590 ;
        RECT 86.575 94.390 136.225 94.590 ;
        RECT 136.575 94.390 152.225 94.590 ;
        RECT 152.575 94.390 154.225 94.590 ;
        RECT 6.890 93.990 7.290 94.390 ;
        RECT 8.890 93.990 9.290 94.390 ;
        RECT 10.890 93.990 11.290 94.390 ;
        RECT 12.890 93.990 13.290 94.390 ;
        RECT 14.890 93.990 15.290 94.390 ;
        RECT 16.890 93.990 17.290 94.390 ;
        RECT 18.890 93.990 19.290 94.390 ;
        RECT 20.890 93.990 21.290 94.390 ;
        RECT 22.890 93.990 23.290 94.390 ;
        RECT 24.890 93.990 25.290 94.390 ;
        RECT 26.890 93.990 27.290 94.390 ;
        RECT 28.890 93.990 29.290 94.390 ;
        RECT 30.890 93.990 31.290 94.390 ;
        RECT 32.890 93.990 33.290 94.390 ;
        RECT 34.890 93.990 35.290 94.390 ;
        RECT 36.890 93.990 37.290 94.390 ;
        RECT 38.890 93.990 39.290 94.390 ;
        RECT 40.890 93.990 41.290 94.390 ;
        RECT 42.890 93.990 43.290 94.390 ;
        RECT 44.890 93.990 45.290 94.390 ;
        RECT 46.890 93.990 47.290 94.390 ;
        RECT 48.890 93.990 49.290 94.390 ;
        RECT 50.890 93.990 51.290 94.390 ;
        RECT 52.890 93.990 53.290 94.390 ;
        RECT 54.890 93.990 55.290 94.390 ;
        RECT 56.890 93.990 57.290 94.390 ;
        RECT 58.890 93.990 59.290 94.390 ;
        RECT 60.890 93.990 61.290 94.390 ;
        RECT 62.890 93.990 63.290 94.390 ;
        RECT 64.890 93.990 65.290 94.390 ;
        RECT 66.890 93.990 67.290 94.390 ;
        RECT 68.890 93.990 69.290 94.390 ;
        RECT 70.890 93.990 71.290 94.390 ;
        RECT 72.890 93.990 73.290 94.390 ;
        RECT 87.825 93.990 88.225 94.390 ;
        RECT 89.825 93.990 90.225 94.390 ;
        RECT 91.825 93.990 92.225 94.390 ;
        RECT 93.825 93.990 94.225 94.390 ;
        RECT 95.825 93.990 96.225 94.390 ;
        RECT 97.825 93.990 98.225 94.390 ;
        RECT 99.825 93.990 100.225 94.390 ;
        RECT 101.825 93.990 102.225 94.390 ;
        RECT 103.825 93.990 104.225 94.390 ;
        RECT 105.825 93.990 106.225 94.390 ;
        RECT 107.825 93.990 108.225 94.390 ;
        RECT 109.825 93.990 110.225 94.390 ;
        RECT 111.825 93.990 112.225 94.390 ;
        RECT 113.825 93.990 114.225 94.390 ;
        RECT 115.825 93.990 116.225 94.390 ;
        RECT 117.825 93.990 118.225 94.390 ;
        RECT 119.825 93.990 120.225 94.390 ;
        RECT 121.825 93.990 122.225 94.390 ;
        RECT 123.825 93.990 124.225 94.390 ;
        RECT 125.825 93.990 126.225 94.390 ;
        RECT 127.825 93.990 128.225 94.390 ;
        RECT 129.825 93.990 130.225 94.390 ;
        RECT 131.825 93.990 132.225 94.390 ;
        RECT 133.825 93.990 134.225 94.390 ;
        RECT 135.825 93.990 136.225 94.390 ;
        RECT 137.825 93.990 138.225 94.390 ;
        RECT 139.825 93.990 140.225 94.390 ;
        RECT 141.825 93.990 142.225 94.390 ;
        RECT 143.825 93.990 144.225 94.390 ;
        RECT 145.825 93.990 146.225 94.390 ;
        RECT 147.825 93.990 148.225 94.390 ;
        RECT 149.825 93.990 150.225 94.390 ;
        RECT 151.825 93.990 152.225 94.390 ;
        RECT 153.825 93.990 154.225 94.390 ;
        RECT 6.960 93.140 7.220 93.990 ;
        RECT 8.990 93.140 9.190 93.990 ;
        RECT 10.990 93.140 11.190 93.990 ;
        RECT 12.990 93.140 13.190 93.990 ;
        RECT 14.990 93.140 15.190 93.990 ;
        RECT 16.990 93.140 17.190 93.990 ;
        RECT 18.990 93.140 19.190 93.990 ;
        RECT 20.990 93.140 21.190 93.990 ;
        RECT 22.990 93.140 23.190 93.990 ;
        RECT 24.990 93.140 25.190 93.990 ;
        RECT 26.990 93.140 27.190 93.990 ;
        RECT 28.990 93.140 29.190 93.990 ;
        RECT 30.990 93.140 31.190 93.990 ;
        RECT 32.990 93.140 33.190 93.990 ;
        RECT 34.990 93.140 35.190 93.990 ;
        RECT 36.990 93.140 37.190 93.990 ;
        RECT 123.925 93.140 124.125 93.990 ;
        RECT 125.925 93.140 126.125 93.990 ;
        RECT 127.925 93.140 128.125 93.990 ;
        RECT 129.925 93.140 130.125 93.990 ;
        RECT 131.925 93.140 132.125 93.990 ;
        RECT 133.925 93.140 134.125 93.990 ;
        RECT 135.925 93.140 136.125 93.990 ;
        RECT 137.925 93.140 138.125 93.990 ;
        RECT 139.925 93.140 140.125 93.990 ;
        RECT 141.925 93.140 142.125 93.990 ;
        RECT 143.925 93.140 144.125 93.990 ;
        RECT 145.925 93.140 146.125 93.990 ;
        RECT 147.925 93.140 148.125 93.990 ;
        RECT 149.925 93.140 150.125 93.990 ;
        RECT 151.925 93.140 152.125 93.990 ;
        RECT 153.895 93.140 154.155 93.990 ;
        RECT 6.890 92.740 7.290 93.140 ;
        RECT 8.890 92.740 9.290 93.140 ;
        RECT 10.890 92.740 11.290 93.140 ;
        RECT 12.890 92.740 13.290 93.140 ;
        RECT 14.890 92.740 15.290 93.140 ;
        RECT 16.890 92.740 17.290 93.140 ;
        RECT 18.890 92.740 19.290 93.140 ;
        RECT 20.890 92.740 21.290 93.140 ;
        RECT 22.890 92.740 23.290 93.140 ;
        RECT 24.890 92.740 25.290 93.140 ;
        RECT 26.890 92.740 27.290 93.140 ;
        RECT 28.890 92.740 29.290 93.140 ;
        RECT 30.890 92.740 31.290 93.140 ;
        RECT 32.890 92.740 33.290 93.140 ;
        RECT 34.890 92.740 35.290 93.140 ;
        RECT 36.890 92.740 37.290 93.140 ;
        RECT 38.890 92.740 39.290 93.140 ;
        RECT 40.890 92.740 41.290 93.140 ;
        RECT 42.890 92.740 43.290 93.140 ;
        RECT 44.890 92.740 45.290 93.140 ;
        RECT 46.890 92.740 47.290 93.140 ;
        RECT 48.890 92.740 49.290 93.140 ;
        RECT 50.890 92.740 51.290 93.140 ;
        RECT 52.890 92.740 53.290 93.140 ;
        RECT 54.890 92.740 55.290 93.140 ;
        RECT 56.890 92.740 57.290 93.140 ;
        RECT 58.890 92.740 59.290 93.140 ;
        RECT 60.890 92.740 61.290 93.140 ;
        RECT 62.890 92.740 63.290 93.140 ;
        RECT 64.890 92.740 65.290 93.140 ;
        RECT 66.890 92.740 67.290 93.140 ;
        RECT 68.890 92.740 69.290 93.140 ;
        RECT 70.890 92.740 71.290 93.140 ;
        RECT 72.890 92.740 73.290 93.140 ;
        RECT 87.825 92.740 88.225 93.140 ;
        RECT 89.825 92.740 90.225 93.140 ;
        RECT 91.825 92.740 92.225 93.140 ;
        RECT 93.825 92.740 94.225 93.140 ;
        RECT 95.825 92.740 96.225 93.140 ;
        RECT 97.825 92.740 98.225 93.140 ;
        RECT 99.825 92.740 100.225 93.140 ;
        RECT 101.825 92.740 102.225 93.140 ;
        RECT 103.825 92.740 104.225 93.140 ;
        RECT 105.825 92.740 106.225 93.140 ;
        RECT 107.825 92.740 108.225 93.140 ;
        RECT 109.825 92.740 110.225 93.140 ;
        RECT 111.825 92.740 112.225 93.140 ;
        RECT 113.825 92.740 114.225 93.140 ;
        RECT 115.825 92.740 116.225 93.140 ;
        RECT 117.825 92.740 118.225 93.140 ;
        RECT 119.825 92.740 120.225 93.140 ;
        RECT 121.825 92.740 122.225 93.140 ;
        RECT 123.825 92.740 124.225 93.140 ;
        RECT 125.825 92.740 126.225 93.140 ;
        RECT 127.825 92.740 128.225 93.140 ;
        RECT 129.825 92.740 130.225 93.140 ;
        RECT 131.825 92.740 132.225 93.140 ;
        RECT 133.825 92.740 134.225 93.140 ;
        RECT 135.825 92.740 136.225 93.140 ;
        RECT 137.825 92.740 138.225 93.140 ;
        RECT 139.825 92.740 140.225 93.140 ;
        RECT 141.825 92.740 142.225 93.140 ;
        RECT 143.825 92.740 144.225 93.140 ;
        RECT 145.825 92.740 146.225 93.140 ;
        RECT 147.825 92.740 148.225 93.140 ;
        RECT 149.825 92.740 150.225 93.140 ;
        RECT 151.825 92.740 152.225 93.140 ;
        RECT 153.825 92.740 154.225 93.140 ;
        RECT 6.890 92.540 8.540 92.740 ;
        RECT 8.890 92.540 24.540 92.740 ;
        RECT 24.890 92.540 38.540 92.740 ;
        RECT 38.890 92.540 74.540 92.740 ;
        RECT 86.575 92.540 122.225 92.740 ;
        RECT 122.575 92.540 136.225 92.740 ;
        RECT 136.575 92.540 152.225 92.740 ;
        RECT 152.575 92.540 154.225 92.740 ;
        RECT 6.890 92.140 7.290 92.540 ;
        RECT 8.890 92.140 9.290 92.540 ;
        RECT 10.890 92.140 11.290 92.540 ;
        RECT 12.890 92.140 13.290 92.540 ;
        RECT 14.890 92.140 15.290 92.540 ;
        RECT 16.890 92.140 17.290 92.540 ;
        RECT 18.890 92.140 19.290 92.540 ;
        RECT 20.890 92.140 21.290 92.540 ;
        RECT 22.890 92.140 23.290 92.540 ;
        RECT 24.890 92.140 25.290 92.540 ;
        RECT 26.890 92.140 27.290 92.540 ;
        RECT 28.890 92.140 29.290 92.540 ;
        RECT 30.890 92.140 31.290 92.540 ;
        RECT 32.890 92.140 33.290 92.540 ;
        RECT 34.890 92.140 35.290 92.540 ;
        RECT 36.890 92.140 37.290 92.540 ;
        RECT 38.890 92.140 39.290 92.540 ;
        RECT 40.890 92.140 41.290 92.540 ;
        RECT 42.890 92.140 43.290 92.540 ;
        RECT 44.890 92.140 45.290 92.540 ;
        RECT 46.890 92.140 47.290 92.540 ;
        RECT 48.890 92.140 49.290 92.540 ;
        RECT 50.890 92.140 51.290 92.540 ;
        RECT 52.890 92.140 53.290 92.540 ;
        RECT 54.890 92.140 55.290 92.540 ;
        RECT 56.890 92.140 57.290 92.540 ;
        RECT 58.890 92.140 59.290 92.540 ;
        RECT 60.890 92.140 61.290 92.540 ;
        RECT 62.890 92.140 63.290 92.540 ;
        RECT 64.890 92.140 65.290 92.540 ;
        RECT 66.890 92.140 67.290 92.540 ;
        RECT 68.890 92.140 69.290 92.540 ;
        RECT 70.890 92.140 71.290 92.540 ;
        RECT 72.890 92.140 73.290 92.540 ;
        RECT 87.825 92.140 88.225 92.540 ;
        RECT 89.825 92.140 90.225 92.540 ;
        RECT 91.825 92.140 92.225 92.540 ;
        RECT 93.825 92.140 94.225 92.540 ;
        RECT 95.825 92.140 96.225 92.540 ;
        RECT 97.825 92.140 98.225 92.540 ;
        RECT 99.825 92.140 100.225 92.540 ;
        RECT 101.825 92.140 102.225 92.540 ;
        RECT 103.825 92.140 104.225 92.540 ;
        RECT 105.825 92.140 106.225 92.540 ;
        RECT 107.825 92.140 108.225 92.540 ;
        RECT 109.825 92.140 110.225 92.540 ;
        RECT 111.825 92.140 112.225 92.540 ;
        RECT 113.825 92.140 114.225 92.540 ;
        RECT 115.825 92.140 116.225 92.540 ;
        RECT 117.825 92.140 118.225 92.540 ;
        RECT 119.825 92.140 120.225 92.540 ;
        RECT 121.825 92.140 122.225 92.540 ;
        RECT 123.825 92.140 124.225 92.540 ;
        RECT 125.825 92.140 126.225 92.540 ;
        RECT 127.825 92.140 128.225 92.540 ;
        RECT 129.825 92.140 130.225 92.540 ;
        RECT 131.825 92.140 132.225 92.540 ;
        RECT 133.825 92.140 134.225 92.540 ;
        RECT 135.825 92.140 136.225 92.540 ;
        RECT 137.825 92.140 138.225 92.540 ;
        RECT 139.825 92.140 140.225 92.540 ;
        RECT 141.825 92.140 142.225 92.540 ;
        RECT 143.825 92.140 144.225 92.540 ;
        RECT 145.825 92.140 146.225 92.540 ;
        RECT 147.825 92.140 148.225 92.540 ;
        RECT 149.825 92.140 150.225 92.540 ;
        RECT 151.825 92.140 152.225 92.540 ;
        RECT 153.825 92.140 154.225 92.540 ;
        RECT 6.960 91.290 7.220 92.140 ;
        RECT 8.990 91.290 9.190 92.140 ;
        RECT 10.990 91.290 11.190 92.140 ;
        RECT 12.990 91.290 13.190 92.140 ;
        RECT 14.990 91.290 15.190 92.140 ;
        RECT 16.990 91.290 17.190 92.140 ;
        RECT 18.990 91.290 19.190 92.140 ;
        RECT 20.990 91.290 21.190 92.140 ;
        RECT 22.990 91.290 23.190 92.140 ;
        RECT 24.990 91.290 25.190 92.140 ;
        RECT 26.990 91.290 27.190 92.140 ;
        RECT 28.990 91.290 29.190 92.140 ;
        RECT 30.990 91.290 31.190 92.140 ;
        RECT 32.990 91.290 33.190 92.140 ;
        RECT 34.990 91.290 35.190 92.140 ;
        RECT 36.990 91.290 37.190 92.140 ;
        RECT 38.990 91.290 39.190 92.140 ;
        RECT 40.990 91.290 41.190 92.140 ;
        RECT 42.990 91.290 43.190 92.140 ;
        RECT 44.990 91.290 45.190 92.140 ;
        RECT 46.990 91.290 47.190 92.140 ;
        RECT 48.990 91.290 49.190 92.140 ;
        RECT 50.990 91.290 51.190 92.140 ;
        RECT 52.990 91.290 53.190 92.140 ;
        RECT 54.990 91.290 55.190 92.140 ;
        RECT 56.990 91.290 57.190 92.140 ;
        RECT 58.990 91.290 59.190 92.140 ;
        RECT 60.990 91.290 61.190 92.140 ;
        RECT 62.990 91.290 63.190 92.140 ;
        RECT 64.990 91.290 65.190 92.140 ;
        RECT 66.990 91.290 67.190 92.140 ;
        RECT 68.990 91.290 69.190 92.140 ;
        RECT 70.990 91.290 71.190 92.140 ;
        RECT 89.925 91.290 90.125 92.140 ;
        RECT 91.925 91.290 92.125 92.140 ;
        RECT 93.925 91.290 94.125 92.140 ;
        RECT 95.925 91.290 96.125 92.140 ;
        RECT 97.925 91.290 98.125 92.140 ;
        RECT 99.925 91.290 100.125 92.140 ;
        RECT 101.925 91.290 102.125 92.140 ;
        RECT 103.925 91.290 104.125 92.140 ;
        RECT 105.925 91.290 106.125 92.140 ;
        RECT 107.925 91.290 108.125 92.140 ;
        RECT 109.925 91.290 110.125 92.140 ;
        RECT 111.925 91.290 112.125 92.140 ;
        RECT 113.925 91.290 114.125 92.140 ;
        RECT 115.925 91.290 116.125 92.140 ;
        RECT 117.925 91.290 118.125 92.140 ;
        RECT 119.925 91.290 120.125 92.140 ;
        RECT 121.925 91.290 122.125 92.140 ;
        RECT 123.925 91.290 124.125 92.140 ;
        RECT 125.925 91.290 126.125 92.140 ;
        RECT 127.925 91.290 128.125 92.140 ;
        RECT 129.925 91.290 130.125 92.140 ;
        RECT 131.925 91.290 132.125 92.140 ;
        RECT 133.925 91.290 134.125 92.140 ;
        RECT 135.925 91.290 136.125 92.140 ;
        RECT 137.925 91.290 138.125 92.140 ;
        RECT 139.925 91.290 140.125 92.140 ;
        RECT 141.925 91.290 142.125 92.140 ;
        RECT 143.925 91.290 144.125 92.140 ;
        RECT 145.925 91.290 146.125 92.140 ;
        RECT 147.925 91.290 148.125 92.140 ;
        RECT 149.925 91.290 150.125 92.140 ;
        RECT 151.925 91.290 152.125 92.140 ;
        RECT 153.895 91.290 154.155 92.140 ;
        RECT 6.890 90.890 7.290 91.290 ;
        RECT 8.890 90.890 9.290 91.290 ;
        RECT 10.890 90.890 11.290 91.290 ;
        RECT 12.890 90.890 13.290 91.290 ;
        RECT 14.890 90.890 15.290 91.290 ;
        RECT 16.890 90.890 17.290 91.290 ;
        RECT 18.890 90.890 19.290 91.290 ;
        RECT 20.890 90.890 21.290 91.290 ;
        RECT 22.890 90.890 23.290 91.290 ;
        RECT 24.890 90.890 25.290 91.290 ;
        RECT 26.890 90.890 27.290 91.290 ;
        RECT 28.890 90.890 29.290 91.290 ;
        RECT 30.890 90.890 31.290 91.290 ;
        RECT 32.890 90.890 33.290 91.290 ;
        RECT 34.890 90.890 35.290 91.290 ;
        RECT 36.890 90.890 37.290 91.290 ;
        RECT 38.890 90.890 39.290 91.290 ;
        RECT 40.890 90.890 41.290 91.290 ;
        RECT 42.890 90.890 43.290 91.290 ;
        RECT 44.890 90.890 45.290 91.290 ;
        RECT 46.890 90.890 47.290 91.290 ;
        RECT 48.890 90.890 49.290 91.290 ;
        RECT 50.890 90.890 51.290 91.290 ;
        RECT 52.890 90.890 53.290 91.290 ;
        RECT 54.890 90.890 55.290 91.290 ;
        RECT 56.890 90.890 57.290 91.290 ;
        RECT 58.890 90.890 59.290 91.290 ;
        RECT 60.890 90.890 61.290 91.290 ;
        RECT 62.890 90.890 63.290 91.290 ;
        RECT 64.890 90.890 65.290 91.290 ;
        RECT 66.890 90.890 67.290 91.290 ;
        RECT 68.890 90.890 69.290 91.290 ;
        RECT 70.890 90.890 71.290 91.290 ;
        RECT 72.890 90.890 73.290 91.290 ;
        RECT 87.825 90.890 88.225 91.290 ;
        RECT 89.825 90.890 90.225 91.290 ;
        RECT 91.825 90.890 92.225 91.290 ;
        RECT 93.825 90.890 94.225 91.290 ;
        RECT 95.825 90.890 96.225 91.290 ;
        RECT 97.825 90.890 98.225 91.290 ;
        RECT 99.825 90.890 100.225 91.290 ;
        RECT 101.825 90.890 102.225 91.290 ;
        RECT 103.825 90.890 104.225 91.290 ;
        RECT 105.825 90.890 106.225 91.290 ;
        RECT 107.825 90.890 108.225 91.290 ;
        RECT 109.825 90.890 110.225 91.290 ;
        RECT 111.825 90.890 112.225 91.290 ;
        RECT 113.825 90.890 114.225 91.290 ;
        RECT 115.825 90.890 116.225 91.290 ;
        RECT 117.825 90.890 118.225 91.290 ;
        RECT 119.825 90.890 120.225 91.290 ;
        RECT 121.825 90.890 122.225 91.290 ;
        RECT 123.825 90.890 124.225 91.290 ;
        RECT 125.825 90.890 126.225 91.290 ;
        RECT 127.825 90.890 128.225 91.290 ;
        RECT 129.825 90.890 130.225 91.290 ;
        RECT 131.825 90.890 132.225 91.290 ;
        RECT 133.825 90.890 134.225 91.290 ;
        RECT 135.825 90.890 136.225 91.290 ;
        RECT 137.825 90.890 138.225 91.290 ;
        RECT 139.825 90.890 140.225 91.290 ;
        RECT 141.825 90.890 142.225 91.290 ;
        RECT 143.825 90.890 144.225 91.290 ;
        RECT 145.825 90.890 146.225 91.290 ;
        RECT 147.825 90.890 148.225 91.290 ;
        RECT 149.825 90.890 150.225 91.290 ;
        RECT 151.825 90.890 152.225 91.290 ;
        RECT 153.825 90.890 154.225 91.290 ;
        RECT 6.890 90.690 8.540 90.890 ;
        RECT 8.890 90.690 24.540 90.890 ;
        RECT 24.890 90.690 38.540 90.890 ;
        RECT 38.890 90.690 74.540 90.890 ;
        RECT 86.575 90.690 122.225 90.890 ;
        RECT 122.575 90.690 136.225 90.890 ;
        RECT 136.575 90.690 152.225 90.890 ;
        RECT 152.575 90.690 154.225 90.890 ;
        RECT 6.890 90.290 7.290 90.690 ;
        RECT 8.890 90.290 9.290 90.690 ;
        RECT 10.890 90.290 11.290 90.690 ;
        RECT 12.890 90.290 13.290 90.690 ;
        RECT 14.890 90.290 15.290 90.690 ;
        RECT 16.890 90.290 17.290 90.690 ;
        RECT 18.890 90.290 19.290 90.690 ;
        RECT 20.890 90.290 21.290 90.690 ;
        RECT 22.890 90.290 23.290 90.690 ;
        RECT 24.890 90.290 25.290 90.690 ;
        RECT 26.890 90.290 27.290 90.690 ;
        RECT 28.890 90.290 29.290 90.690 ;
        RECT 30.890 90.290 31.290 90.690 ;
        RECT 32.890 90.290 33.290 90.690 ;
        RECT 34.890 90.290 35.290 90.690 ;
        RECT 36.890 90.290 37.290 90.690 ;
        RECT 38.890 90.290 39.290 90.690 ;
        RECT 40.890 90.290 41.290 90.690 ;
        RECT 42.890 90.290 43.290 90.690 ;
        RECT 44.890 90.290 45.290 90.690 ;
        RECT 46.890 90.290 47.290 90.690 ;
        RECT 48.890 90.290 49.290 90.690 ;
        RECT 50.890 90.290 51.290 90.690 ;
        RECT 52.890 90.290 53.290 90.690 ;
        RECT 54.890 90.290 55.290 90.690 ;
        RECT 56.890 90.290 57.290 90.690 ;
        RECT 58.890 90.290 59.290 90.690 ;
        RECT 60.890 90.290 61.290 90.690 ;
        RECT 62.890 90.290 63.290 90.690 ;
        RECT 64.890 90.290 65.290 90.690 ;
        RECT 66.890 90.290 67.290 90.690 ;
        RECT 68.890 90.290 69.290 90.690 ;
        RECT 70.890 90.290 71.290 90.690 ;
        RECT 72.890 90.290 73.290 90.690 ;
        RECT 87.825 90.290 88.225 90.690 ;
        RECT 89.825 90.290 90.225 90.690 ;
        RECT 91.825 90.290 92.225 90.690 ;
        RECT 93.825 90.290 94.225 90.690 ;
        RECT 95.825 90.290 96.225 90.690 ;
        RECT 97.825 90.290 98.225 90.690 ;
        RECT 99.825 90.290 100.225 90.690 ;
        RECT 101.825 90.290 102.225 90.690 ;
        RECT 103.825 90.290 104.225 90.690 ;
        RECT 105.825 90.290 106.225 90.690 ;
        RECT 107.825 90.290 108.225 90.690 ;
        RECT 109.825 90.290 110.225 90.690 ;
        RECT 111.825 90.290 112.225 90.690 ;
        RECT 113.825 90.290 114.225 90.690 ;
        RECT 115.825 90.290 116.225 90.690 ;
        RECT 117.825 90.290 118.225 90.690 ;
        RECT 119.825 90.290 120.225 90.690 ;
        RECT 121.825 90.290 122.225 90.690 ;
        RECT 123.825 90.290 124.225 90.690 ;
        RECT 125.825 90.290 126.225 90.690 ;
        RECT 127.825 90.290 128.225 90.690 ;
        RECT 129.825 90.290 130.225 90.690 ;
        RECT 131.825 90.290 132.225 90.690 ;
        RECT 133.825 90.290 134.225 90.690 ;
        RECT 135.825 90.290 136.225 90.690 ;
        RECT 137.825 90.290 138.225 90.690 ;
        RECT 139.825 90.290 140.225 90.690 ;
        RECT 141.825 90.290 142.225 90.690 ;
        RECT 143.825 90.290 144.225 90.690 ;
        RECT 145.825 90.290 146.225 90.690 ;
        RECT 147.825 90.290 148.225 90.690 ;
        RECT 149.825 90.290 150.225 90.690 ;
        RECT 151.825 90.290 152.225 90.690 ;
        RECT 153.825 90.290 154.225 90.690 ;
        RECT 6.960 89.440 7.220 90.290 ;
        RECT 8.990 89.440 9.190 90.290 ;
        RECT 10.990 89.440 11.190 90.290 ;
        RECT 12.990 89.440 13.190 90.290 ;
        RECT 14.990 89.440 15.190 90.290 ;
        RECT 16.990 89.440 17.190 90.290 ;
        RECT 18.990 89.440 19.190 90.290 ;
        RECT 20.990 89.440 21.190 90.290 ;
        RECT 22.990 89.440 23.190 90.290 ;
        RECT 24.990 89.440 25.190 90.290 ;
        RECT 26.990 89.440 27.190 90.290 ;
        RECT 28.990 89.440 29.190 90.290 ;
        RECT 30.990 89.440 31.190 90.290 ;
        RECT 32.990 89.440 33.190 90.290 ;
        RECT 34.990 89.440 35.190 90.290 ;
        RECT 36.990 89.440 37.190 90.290 ;
        RECT 38.990 89.440 39.190 90.290 ;
        RECT 40.990 89.440 41.190 90.290 ;
        RECT 42.990 89.440 43.190 90.290 ;
        RECT 44.990 89.440 45.190 90.290 ;
        RECT 46.990 89.440 47.190 90.290 ;
        RECT 48.990 89.440 49.190 90.290 ;
        RECT 50.990 89.440 51.190 90.290 ;
        RECT 52.990 89.440 53.190 90.290 ;
        RECT 54.990 89.440 55.190 90.290 ;
        RECT 56.990 89.440 57.190 90.290 ;
        RECT 58.990 89.440 59.190 90.290 ;
        RECT 60.990 89.440 61.190 90.290 ;
        RECT 62.990 89.440 63.190 90.290 ;
        RECT 64.990 89.440 65.190 90.290 ;
        RECT 66.990 89.440 67.190 90.290 ;
        RECT 68.990 89.440 69.190 90.290 ;
        RECT 70.990 89.440 71.190 90.290 ;
        RECT 89.925 89.440 90.125 90.290 ;
        RECT 91.925 89.440 92.125 90.290 ;
        RECT 93.925 89.440 94.125 90.290 ;
        RECT 95.925 89.440 96.125 90.290 ;
        RECT 97.925 89.440 98.125 90.290 ;
        RECT 99.925 89.440 100.125 90.290 ;
        RECT 101.925 89.440 102.125 90.290 ;
        RECT 103.925 89.440 104.125 90.290 ;
        RECT 105.925 89.440 106.125 90.290 ;
        RECT 107.925 89.440 108.125 90.290 ;
        RECT 109.925 89.440 110.125 90.290 ;
        RECT 111.925 89.440 112.125 90.290 ;
        RECT 113.925 89.440 114.125 90.290 ;
        RECT 115.925 89.440 116.125 90.290 ;
        RECT 117.925 89.440 118.125 90.290 ;
        RECT 119.925 89.440 120.125 90.290 ;
        RECT 121.925 89.440 122.125 90.290 ;
        RECT 123.925 89.440 124.125 90.290 ;
        RECT 125.925 89.440 126.125 90.290 ;
        RECT 127.925 89.440 128.125 90.290 ;
        RECT 129.925 89.440 130.125 90.290 ;
        RECT 131.925 89.440 132.125 90.290 ;
        RECT 133.925 89.440 134.125 90.290 ;
        RECT 135.925 89.440 136.125 90.290 ;
        RECT 137.925 89.440 138.125 90.290 ;
        RECT 139.925 89.440 140.125 90.290 ;
        RECT 141.925 89.440 142.125 90.290 ;
        RECT 143.925 89.440 144.125 90.290 ;
        RECT 145.925 89.440 146.125 90.290 ;
        RECT 147.925 89.440 148.125 90.290 ;
        RECT 149.925 89.440 150.125 90.290 ;
        RECT 151.925 89.440 152.125 90.290 ;
        RECT 153.895 89.440 154.155 90.290 ;
        RECT 6.890 89.040 7.290 89.440 ;
        RECT 8.890 89.040 9.290 89.440 ;
        RECT 10.890 89.040 11.290 89.440 ;
        RECT 12.890 89.040 13.290 89.440 ;
        RECT 14.890 89.040 15.290 89.440 ;
        RECT 16.890 89.040 17.290 89.440 ;
        RECT 18.890 89.040 19.290 89.440 ;
        RECT 20.890 89.040 21.290 89.440 ;
        RECT 22.890 89.040 23.290 89.440 ;
        RECT 24.890 89.040 25.290 89.440 ;
        RECT 26.890 89.040 27.290 89.440 ;
        RECT 28.890 89.040 29.290 89.440 ;
        RECT 30.890 89.040 31.290 89.440 ;
        RECT 32.890 89.040 33.290 89.440 ;
        RECT 34.890 89.040 35.290 89.440 ;
        RECT 36.890 89.040 37.290 89.440 ;
        RECT 38.890 89.040 39.290 89.440 ;
        RECT 40.890 89.040 41.290 89.440 ;
        RECT 42.890 89.040 43.290 89.440 ;
        RECT 44.890 89.040 45.290 89.440 ;
        RECT 46.890 89.040 47.290 89.440 ;
        RECT 48.890 89.040 49.290 89.440 ;
        RECT 50.890 89.040 51.290 89.440 ;
        RECT 52.890 89.040 53.290 89.440 ;
        RECT 54.890 89.040 55.290 89.440 ;
        RECT 56.890 89.040 57.290 89.440 ;
        RECT 58.890 89.040 59.290 89.440 ;
        RECT 60.890 89.040 61.290 89.440 ;
        RECT 62.890 89.040 63.290 89.440 ;
        RECT 64.890 89.040 65.290 89.440 ;
        RECT 66.890 89.040 67.290 89.440 ;
        RECT 68.890 89.040 69.290 89.440 ;
        RECT 70.890 89.040 71.290 89.440 ;
        RECT 72.890 89.040 73.290 89.440 ;
        RECT 87.825 89.040 88.225 89.440 ;
        RECT 89.825 89.040 90.225 89.440 ;
        RECT 91.825 89.040 92.225 89.440 ;
        RECT 93.825 89.040 94.225 89.440 ;
        RECT 95.825 89.040 96.225 89.440 ;
        RECT 97.825 89.040 98.225 89.440 ;
        RECT 99.825 89.040 100.225 89.440 ;
        RECT 101.825 89.040 102.225 89.440 ;
        RECT 103.825 89.040 104.225 89.440 ;
        RECT 105.825 89.040 106.225 89.440 ;
        RECT 107.825 89.040 108.225 89.440 ;
        RECT 109.825 89.040 110.225 89.440 ;
        RECT 111.825 89.040 112.225 89.440 ;
        RECT 113.825 89.040 114.225 89.440 ;
        RECT 115.825 89.040 116.225 89.440 ;
        RECT 117.825 89.040 118.225 89.440 ;
        RECT 119.825 89.040 120.225 89.440 ;
        RECT 121.825 89.040 122.225 89.440 ;
        RECT 123.825 89.040 124.225 89.440 ;
        RECT 125.825 89.040 126.225 89.440 ;
        RECT 127.825 89.040 128.225 89.440 ;
        RECT 129.825 89.040 130.225 89.440 ;
        RECT 131.825 89.040 132.225 89.440 ;
        RECT 133.825 89.040 134.225 89.440 ;
        RECT 135.825 89.040 136.225 89.440 ;
        RECT 137.825 89.040 138.225 89.440 ;
        RECT 139.825 89.040 140.225 89.440 ;
        RECT 141.825 89.040 142.225 89.440 ;
        RECT 143.825 89.040 144.225 89.440 ;
        RECT 145.825 89.040 146.225 89.440 ;
        RECT 147.825 89.040 148.225 89.440 ;
        RECT 149.825 89.040 150.225 89.440 ;
        RECT 151.825 89.040 152.225 89.440 ;
        RECT 153.825 89.040 154.225 89.440 ;
        RECT 6.890 88.840 8.540 89.040 ;
        RECT 8.890 88.840 24.540 89.040 ;
        RECT 24.890 88.840 38.540 89.040 ;
        RECT 38.890 88.840 74.540 89.040 ;
        RECT 86.575 88.840 122.225 89.040 ;
        RECT 122.575 88.840 136.225 89.040 ;
        RECT 136.575 88.840 152.225 89.040 ;
        RECT 152.575 88.840 154.225 89.040 ;
        RECT 6.890 88.440 7.290 88.840 ;
        RECT 8.890 88.440 9.290 88.840 ;
        RECT 10.890 88.440 11.290 88.840 ;
        RECT 12.890 88.440 13.290 88.840 ;
        RECT 14.890 88.440 15.290 88.840 ;
        RECT 16.890 88.440 17.290 88.840 ;
        RECT 18.890 88.440 19.290 88.840 ;
        RECT 20.890 88.440 21.290 88.840 ;
        RECT 22.890 88.440 23.290 88.840 ;
        RECT 24.890 88.440 25.290 88.840 ;
        RECT 26.890 88.440 27.290 88.840 ;
        RECT 28.890 88.440 29.290 88.840 ;
        RECT 30.890 88.440 31.290 88.840 ;
        RECT 32.890 88.440 33.290 88.840 ;
        RECT 34.890 88.440 35.290 88.840 ;
        RECT 36.890 88.440 37.290 88.840 ;
        RECT 38.890 88.440 39.290 88.840 ;
        RECT 40.890 88.440 41.290 88.840 ;
        RECT 42.890 88.440 43.290 88.840 ;
        RECT 44.890 88.440 45.290 88.840 ;
        RECT 46.890 88.440 47.290 88.840 ;
        RECT 48.890 88.440 49.290 88.840 ;
        RECT 50.890 88.440 51.290 88.840 ;
        RECT 52.890 88.440 53.290 88.840 ;
        RECT 54.890 88.440 55.290 88.840 ;
        RECT 56.890 88.440 57.290 88.840 ;
        RECT 58.890 88.440 59.290 88.840 ;
        RECT 60.890 88.440 61.290 88.840 ;
        RECT 62.890 88.440 63.290 88.840 ;
        RECT 64.890 88.440 65.290 88.840 ;
        RECT 66.890 88.440 67.290 88.840 ;
        RECT 68.890 88.440 69.290 88.840 ;
        RECT 70.890 88.440 71.290 88.840 ;
        RECT 72.890 88.440 73.290 88.840 ;
        RECT 87.825 88.440 88.225 88.840 ;
        RECT 89.825 88.440 90.225 88.840 ;
        RECT 91.825 88.440 92.225 88.840 ;
        RECT 93.825 88.440 94.225 88.840 ;
        RECT 95.825 88.440 96.225 88.840 ;
        RECT 97.825 88.440 98.225 88.840 ;
        RECT 99.825 88.440 100.225 88.840 ;
        RECT 101.825 88.440 102.225 88.840 ;
        RECT 103.825 88.440 104.225 88.840 ;
        RECT 105.825 88.440 106.225 88.840 ;
        RECT 107.825 88.440 108.225 88.840 ;
        RECT 109.825 88.440 110.225 88.840 ;
        RECT 111.825 88.440 112.225 88.840 ;
        RECT 113.825 88.440 114.225 88.840 ;
        RECT 115.825 88.440 116.225 88.840 ;
        RECT 117.825 88.440 118.225 88.840 ;
        RECT 119.825 88.440 120.225 88.840 ;
        RECT 121.825 88.440 122.225 88.840 ;
        RECT 123.825 88.440 124.225 88.840 ;
        RECT 125.825 88.440 126.225 88.840 ;
        RECT 127.825 88.440 128.225 88.840 ;
        RECT 129.825 88.440 130.225 88.840 ;
        RECT 131.825 88.440 132.225 88.840 ;
        RECT 133.825 88.440 134.225 88.840 ;
        RECT 135.825 88.440 136.225 88.840 ;
        RECT 137.825 88.440 138.225 88.840 ;
        RECT 139.825 88.440 140.225 88.840 ;
        RECT 141.825 88.440 142.225 88.840 ;
        RECT 143.825 88.440 144.225 88.840 ;
        RECT 145.825 88.440 146.225 88.840 ;
        RECT 147.825 88.440 148.225 88.840 ;
        RECT 149.825 88.440 150.225 88.840 ;
        RECT 151.825 88.440 152.225 88.840 ;
        RECT 153.825 88.440 154.225 88.840 ;
        RECT 6.960 87.590 7.220 88.440 ;
        RECT 8.990 87.590 9.190 88.440 ;
        RECT 10.990 87.590 11.190 88.440 ;
        RECT 12.990 87.590 13.190 88.440 ;
        RECT 14.990 87.590 15.190 88.440 ;
        RECT 16.990 87.590 17.190 88.440 ;
        RECT 18.990 87.590 19.190 88.440 ;
        RECT 20.990 87.590 21.190 88.440 ;
        RECT 22.990 87.590 23.190 88.440 ;
        RECT 24.990 87.590 25.190 88.440 ;
        RECT 26.990 87.590 27.190 88.440 ;
        RECT 28.990 87.590 29.190 88.440 ;
        RECT 30.990 87.590 31.190 88.440 ;
        RECT 32.990 87.590 33.190 88.440 ;
        RECT 34.990 87.590 35.190 88.440 ;
        RECT 36.990 87.590 37.190 88.440 ;
        RECT 38.990 87.590 39.190 88.440 ;
        RECT 40.990 87.590 41.190 88.440 ;
        RECT 42.990 87.590 43.190 88.440 ;
        RECT 44.990 87.590 45.190 88.440 ;
        RECT 46.990 87.590 47.190 88.440 ;
        RECT 48.990 87.590 49.190 88.440 ;
        RECT 50.990 87.590 51.190 88.440 ;
        RECT 52.990 87.590 53.190 88.440 ;
        RECT 54.990 87.590 55.190 88.440 ;
        RECT 56.990 87.590 57.190 88.440 ;
        RECT 58.990 87.590 59.190 88.440 ;
        RECT 60.990 87.590 61.190 88.440 ;
        RECT 62.990 87.590 63.190 88.440 ;
        RECT 64.990 87.590 65.190 88.440 ;
        RECT 66.990 87.590 67.190 88.440 ;
        RECT 68.990 87.590 69.190 88.440 ;
        RECT 70.990 87.590 71.190 88.440 ;
        RECT 89.925 87.590 90.125 88.440 ;
        RECT 91.925 87.590 92.125 88.440 ;
        RECT 93.925 87.590 94.125 88.440 ;
        RECT 95.925 87.590 96.125 88.440 ;
        RECT 97.925 87.590 98.125 88.440 ;
        RECT 99.925 87.590 100.125 88.440 ;
        RECT 101.925 87.590 102.125 88.440 ;
        RECT 103.925 87.590 104.125 88.440 ;
        RECT 105.925 87.590 106.125 88.440 ;
        RECT 107.925 87.590 108.125 88.440 ;
        RECT 109.925 87.590 110.125 88.440 ;
        RECT 111.925 87.590 112.125 88.440 ;
        RECT 113.925 87.590 114.125 88.440 ;
        RECT 115.925 87.590 116.125 88.440 ;
        RECT 117.925 87.590 118.125 88.440 ;
        RECT 119.925 87.590 120.125 88.440 ;
        RECT 121.925 87.590 122.125 88.440 ;
        RECT 123.925 87.590 124.125 88.440 ;
        RECT 125.925 87.590 126.125 88.440 ;
        RECT 127.925 87.590 128.125 88.440 ;
        RECT 129.925 87.590 130.125 88.440 ;
        RECT 131.925 87.590 132.125 88.440 ;
        RECT 133.925 87.590 134.125 88.440 ;
        RECT 135.925 87.590 136.125 88.440 ;
        RECT 137.925 87.590 138.125 88.440 ;
        RECT 139.925 87.590 140.125 88.440 ;
        RECT 141.925 87.590 142.125 88.440 ;
        RECT 143.925 87.590 144.125 88.440 ;
        RECT 145.925 87.590 146.125 88.440 ;
        RECT 147.925 87.590 148.125 88.440 ;
        RECT 149.925 87.590 150.125 88.440 ;
        RECT 151.925 87.590 152.125 88.440 ;
        RECT 153.895 87.590 154.155 88.440 ;
        RECT 6.890 87.190 7.290 87.590 ;
        RECT 8.890 87.190 9.290 87.590 ;
        RECT 10.890 87.190 11.290 87.590 ;
        RECT 12.890 87.190 13.290 87.590 ;
        RECT 14.890 87.190 15.290 87.590 ;
        RECT 16.890 87.190 17.290 87.590 ;
        RECT 18.890 87.190 19.290 87.590 ;
        RECT 20.890 87.190 21.290 87.590 ;
        RECT 22.890 87.190 23.290 87.590 ;
        RECT 24.890 87.190 25.290 87.590 ;
        RECT 26.890 87.190 27.290 87.590 ;
        RECT 28.890 87.190 29.290 87.590 ;
        RECT 30.890 87.190 31.290 87.590 ;
        RECT 32.890 87.190 33.290 87.590 ;
        RECT 34.890 87.190 35.290 87.590 ;
        RECT 36.890 87.190 37.290 87.590 ;
        RECT 38.890 87.190 39.290 87.590 ;
        RECT 40.890 87.190 41.290 87.590 ;
        RECT 42.890 87.190 43.290 87.590 ;
        RECT 44.890 87.190 45.290 87.590 ;
        RECT 46.890 87.190 47.290 87.590 ;
        RECT 48.890 87.190 49.290 87.590 ;
        RECT 50.890 87.190 51.290 87.590 ;
        RECT 52.890 87.190 53.290 87.590 ;
        RECT 54.890 87.190 55.290 87.590 ;
        RECT 56.890 87.190 57.290 87.590 ;
        RECT 58.890 87.190 59.290 87.590 ;
        RECT 60.890 87.190 61.290 87.590 ;
        RECT 62.890 87.190 63.290 87.590 ;
        RECT 64.890 87.190 65.290 87.590 ;
        RECT 66.890 87.190 67.290 87.590 ;
        RECT 68.890 87.190 69.290 87.590 ;
        RECT 70.890 87.190 71.290 87.590 ;
        RECT 72.890 87.190 73.290 87.590 ;
        RECT 87.825 87.190 88.225 87.590 ;
        RECT 89.825 87.190 90.225 87.590 ;
        RECT 91.825 87.190 92.225 87.590 ;
        RECT 93.825 87.190 94.225 87.590 ;
        RECT 95.825 87.190 96.225 87.590 ;
        RECT 97.825 87.190 98.225 87.590 ;
        RECT 99.825 87.190 100.225 87.590 ;
        RECT 101.825 87.190 102.225 87.590 ;
        RECT 103.825 87.190 104.225 87.590 ;
        RECT 105.825 87.190 106.225 87.590 ;
        RECT 107.825 87.190 108.225 87.590 ;
        RECT 109.825 87.190 110.225 87.590 ;
        RECT 111.825 87.190 112.225 87.590 ;
        RECT 113.825 87.190 114.225 87.590 ;
        RECT 115.825 87.190 116.225 87.590 ;
        RECT 117.825 87.190 118.225 87.590 ;
        RECT 119.825 87.190 120.225 87.590 ;
        RECT 121.825 87.190 122.225 87.590 ;
        RECT 123.825 87.190 124.225 87.590 ;
        RECT 125.825 87.190 126.225 87.590 ;
        RECT 127.825 87.190 128.225 87.590 ;
        RECT 129.825 87.190 130.225 87.590 ;
        RECT 131.825 87.190 132.225 87.590 ;
        RECT 133.825 87.190 134.225 87.590 ;
        RECT 135.825 87.190 136.225 87.590 ;
        RECT 137.825 87.190 138.225 87.590 ;
        RECT 139.825 87.190 140.225 87.590 ;
        RECT 141.825 87.190 142.225 87.590 ;
        RECT 143.825 87.190 144.225 87.590 ;
        RECT 145.825 87.190 146.225 87.590 ;
        RECT 147.825 87.190 148.225 87.590 ;
        RECT 149.825 87.190 150.225 87.590 ;
        RECT 151.825 87.190 152.225 87.590 ;
        RECT 153.825 87.190 154.225 87.590 ;
        RECT 6.890 86.990 8.540 87.190 ;
        RECT 8.890 86.990 24.540 87.190 ;
        RECT 24.890 86.990 38.540 87.190 ;
        RECT 38.890 86.990 74.540 87.190 ;
        RECT 86.575 86.990 122.225 87.190 ;
        RECT 122.575 86.990 136.225 87.190 ;
        RECT 136.575 86.990 152.225 87.190 ;
        RECT 152.575 86.990 154.225 87.190 ;
        RECT 6.890 86.590 7.290 86.990 ;
        RECT 8.890 86.590 9.290 86.990 ;
        RECT 10.890 86.590 11.290 86.990 ;
        RECT 12.890 86.590 13.290 86.990 ;
        RECT 14.890 86.590 15.290 86.990 ;
        RECT 16.890 86.590 17.290 86.990 ;
        RECT 18.890 86.590 19.290 86.990 ;
        RECT 20.890 86.590 21.290 86.990 ;
        RECT 22.890 86.590 23.290 86.990 ;
        RECT 24.890 86.590 25.290 86.990 ;
        RECT 26.890 86.590 27.290 86.990 ;
        RECT 28.890 86.590 29.290 86.990 ;
        RECT 30.890 86.590 31.290 86.990 ;
        RECT 32.890 86.590 33.290 86.990 ;
        RECT 34.890 86.590 35.290 86.990 ;
        RECT 36.890 86.590 37.290 86.990 ;
        RECT 38.890 86.590 39.290 86.990 ;
        RECT 40.890 86.590 41.290 86.990 ;
        RECT 42.890 86.590 43.290 86.990 ;
        RECT 44.890 86.590 45.290 86.990 ;
        RECT 46.890 86.590 47.290 86.990 ;
        RECT 48.890 86.590 49.290 86.990 ;
        RECT 50.890 86.590 51.290 86.990 ;
        RECT 52.890 86.590 53.290 86.990 ;
        RECT 54.890 86.590 55.290 86.990 ;
        RECT 56.890 86.590 57.290 86.990 ;
        RECT 58.890 86.590 59.290 86.990 ;
        RECT 60.890 86.590 61.290 86.990 ;
        RECT 62.890 86.590 63.290 86.990 ;
        RECT 64.890 86.590 65.290 86.990 ;
        RECT 66.890 86.590 67.290 86.990 ;
        RECT 68.890 86.590 69.290 86.990 ;
        RECT 70.890 86.590 71.290 86.990 ;
        RECT 72.890 86.590 73.290 86.990 ;
        RECT 87.825 86.590 88.225 86.990 ;
        RECT 89.825 86.590 90.225 86.990 ;
        RECT 91.825 86.590 92.225 86.990 ;
        RECT 93.825 86.590 94.225 86.990 ;
        RECT 95.825 86.590 96.225 86.990 ;
        RECT 97.825 86.590 98.225 86.990 ;
        RECT 99.825 86.590 100.225 86.990 ;
        RECT 101.825 86.590 102.225 86.990 ;
        RECT 103.825 86.590 104.225 86.990 ;
        RECT 105.825 86.590 106.225 86.990 ;
        RECT 107.825 86.590 108.225 86.990 ;
        RECT 109.825 86.590 110.225 86.990 ;
        RECT 111.825 86.590 112.225 86.990 ;
        RECT 113.825 86.590 114.225 86.990 ;
        RECT 115.825 86.590 116.225 86.990 ;
        RECT 117.825 86.590 118.225 86.990 ;
        RECT 119.825 86.590 120.225 86.990 ;
        RECT 121.825 86.590 122.225 86.990 ;
        RECT 123.825 86.590 124.225 86.990 ;
        RECT 125.825 86.590 126.225 86.990 ;
        RECT 127.825 86.590 128.225 86.990 ;
        RECT 129.825 86.590 130.225 86.990 ;
        RECT 131.825 86.590 132.225 86.990 ;
        RECT 133.825 86.590 134.225 86.990 ;
        RECT 135.825 86.590 136.225 86.990 ;
        RECT 137.825 86.590 138.225 86.990 ;
        RECT 139.825 86.590 140.225 86.990 ;
        RECT 141.825 86.590 142.225 86.990 ;
        RECT 143.825 86.590 144.225 86.990 ;
        RECT 145.825 86.590 146.225 86.990 ;
        RECT 147.825 86.590 148.225 86.990 ;
        RECT 149.825 86.590 150.225 86.990 ;
        RECT 151.825 86.590 152.225 86.990 ;
        RECT 153.825 86.590 154.225 86.990 ;
        RECT 6.960 85.740 7.220 86.590 ;
        RECT 8.990 85.740 9.190 86.590 ;
        RECT 10.990 85.740 11.190 86.590 ;
        RECT 12.990 85.740 13.190 86.590 ;
        RECT 14.990 85.740 15.190 86.590 ;
        RECT 16.990 85.740 17.190 86.590 ;
        RECT 18.990 85.740 19.190 86.590 ;
        RECT 20.990 85.740 21.190 86.590 ;
        RECT 22.990 85.740 23.190 86.590 ;
        RECT 24.990 85.740 25.190 86.590 ;
        RECT 26.990 85.740 27.190 86.590 ;
        RECT 28.990 85.740 29.190 86.590 ;
        RECT 30.990 85.740 31.190 86.590 ;
        RECT 32.990 85.740 33.190 86.590 ;
        RECT 34.990 85.740 35.190 86.590 ;
        RECT 36.990 85.740 37.190 86.590 ;
        RECT 38.990 85.740 39.190 86.590 ;
        RECT 40.990 85.740 41.190 86.590 ;
        RECT 42.990 85.740 43.190 86.590 ;
        RECT 44.990 85.740 45.190 86.590 ;
        RECT 46.990 85.740 47.190 86.590 ;
        RECT 48.990 85.740 49.190 86.590 ;
        RECT 50.990 85.740 51.190 86.590 ;
        RECT 52.990 85.740 53.190 86.590 ;
        RECT 54.990 85.740 55.190 86.590 ;
        RECT 56.990 85.740 57.190 86.590 ;
        RECT 58.990 85.740 59.190 86.590 ;
        RECT 60.990 85.740 61.190 86.590 ;
        RECT 62.990 85.740 63.190 86.590 ;
        RECT 64.990 85.740 65.190 86.590 ;
        RECT 66.990 85.740 67.190 86.590 ;
        RECT 68.990 85.740 69.190 86.590 ;
        RECT 70.990 85.740 71.190 86.590 ;
        RECT 89.925 85.740 90.125 86.590 ;
        RECT 91.925 85.740 92.125 86.590 ;
        RECT 93.925 85.740 94.125 86.590 ;
        RECT 95.925 85.740 96.125 86.590 ;
        RECT 97.925 85.740 98.125 86.590 ;
        RECT 99.925 85.740 100.125 86.590 ;
        RECT 101.925 85.740 102.125 86.590 ;
        RECT 103.925 85.740 104.125 86.590 ;
        RECT 105.925 85.740 106.125 86.590 ;
        RECT 107.925 85.740 108.125 86.590 ;
        RECT 109.925 85.740 110.125 86.590 ;
        RECT 111.925 85.740 112.125 86.590 ;
        RECT 113.925 85.740 114.125 86.590 ;
        RECT 115.925 85.740 116.125 86.590 ;
        RECT 117.925 85.740 118.125 86.590 ;
        RECT 119.925 85.740 120.125 86.590 ;
        RECT 121.925 85.740 122.125 86.590 ;
        RECT 123.925 85.740 124.125 86.590 ;
        RECT 125.925 85.740 126.125 86.590 ;
        RECT 127.925 85.740 128.125 86.590 ;
        RECT 129.925 85.740 130.125 86.590 ;
        RECT 131.925 85.740 132.125 86.590 ;
        RECT 133.925 85.740 134.125 86.590 ;
        RECT 135.925 85.740 136.125 86.590 ;
        RECT 137.925 85.740 138.125 86.590 ;
        RECT 139.925 85.740 140.125 86.590 ;
        RECT 141.925 85.740 142.125 86.590 ;
        RECT 143.925 85.740 144.125 86.590 ;
        RECT 145.925 85.740 146.125 86.590 ;
        RECT 147.925 85.740 148.125 86.590 ;
        RECT 149.925 85.740 150.125 86.590 ;
        RECT 151.925 85.740 152.125 86.590 ;
        RECT 153.895 85.740 154.155 86.590 ;
        RECT 6.890 85.340 7.290 85.740 ;
        RECT 8.890 85.340 9.290 85.740 ;
        RECT 10.890 85.340 11.290 85.740 ;
        RECT 12.890 85.340 13.290 85.740 ;
        RECT 14.890 85.340 15.290 85.740 ;
        RECT 16.890 85.340 17.290 85.740 ;
        RECT 18.890 85.340 19.290 85.740 ;
        RECT 20.890 85.340 21.290 85.740 ;
        RECT 22.890 85.340 23.290 85.740 ;
        RECT 24.890 85.340 25.290 85.740 ;
        RECT 26.890 85.340 27.290 85.740 ;
        RECT 28.890 85.340 29.290 85.740 ;
        RECT 30.890 85.340 31.290 85.740 ;
        RECT 32.890 85.340 33.290 85.740 ;
        RECT 34.890 85.340 35.290 85.740 ;
        RECT 36.890 85.340 37.290 85.740 ;
        RECT 38.890 85.340 39.290 85.740 ;
        RECT 40.890 85.340 41.290 85.740 ;
        RECT 42.890 85.340 43.290 85.740 ;
        RECT 44.890 85.340 45.290 85.740 ;
        RECT 46.890 85.340 47.290 85.740 ;
        RECT 48.890 85.340 49.290 85.740 ;
        RECT 50.890 85.340 51.290 85.740 ;
        RECT 52.890 85.340 53.290 85.740 ;
        RECT 54.890 85.340 55.290 85.740 ;
        RECT 56.890 85.340 57.290 85.740 ;
        RECT 58.890 85.340 59.290 85.740 ;
        RECT 60.890 85.340 61.290 85.740 ;
        RECT 62.890 85.340 63.290 85.740 ;
        RECT 64.890 85.340 65.290 85.740 ;
        RECT 66.890 85.340 67.290 85.740 ;
        RECT 68.890 85.340 69.290 85.740 ;
        RECT 70.890 85.340 71.290 85.740 ;
        RECT 72.890 85.340 73.290 85.740 ;
        RECT 87.825 85.340 88.225 85.740 ;
        RECT 89.825 85.340 90.225 85.740 ;
        RECT 91.825 85.340 92.225 85.740 ;
        RECT 93.825 85.340 94.225 85.740 ;
        RECT 95.825 85.340 96.225 85.740 ;
        RECT 97.825 85.340 98.225 85.740 ;
        RECT 99.825 85.340 100.225 85.740 ;
        RECT 101.825 85.340 102.225 85.740 ;
        RECT 103.825 85.340 104.225 85.740 ;
        RECT 105.825 85.340 106.225 85.740 ;
        RECT 107.825 85.340 108.225 85.740 ;
        RECT 109.825 85.340 110.225 85.740 ;
        RECT 111.825 85.340 112.225 85.740 ;
        RECT 113.825 85.340 114.225 85.740 ;
        RECT 115.825 85.340 116.225 85.740 ;
        RECT 117.825 85.340 118.225 85.740 ;
        RECT 119.825 85.340 120.225 85.740 ;
        RECT 121.825 85.340 122.225 85.740 ;
        RECT 123.825 85.340 124.225 85.740 ;
        RECT 125.825 85.340 126.225 85.740 ;
        RECT 127.825 85.340 128.225 85.740 ;
        RECT 129.825 85.340 130.225 85.740 ;
        RECT 131.825 85.340 132.225 85.740 ;
        RECT 133.825 85.340 134.225 85.740 ;
        RECT 135.825 85.340 136.225 85.740 ;
        RECT 137.825 85.340 138.225 85.740 ;
        RECT 139.825 85.340 140.225 85.740 ;
        RECT 141.825 85.340 142.225 85.740 ;
        RECT 143.825 85.340 144.225 85.740 ;
        RECT 145.825 85.340 146.225 85.740 ;
        RECT 147.825 85.340 148.225 85.740 ;
        RECT 149.825 85.340 150.225 85.740 ;
        RECT 151.825 85.340 152.225 85.740 ;
        RECT 153.825 85.340 154.225 85.740 ;
        RECT 6.890 85.140 8.540 85.340 ;
        RECT 8.890 85.140 24.540 85.340 ;
        RECT 24.890 85.140 38.540 85.340 ;
        RECT 38.890 85.140 74.540 85.340 ;
        RECT 86.575 85.140 122.225 85.340 ;
        RECT 122.575 85.140 136.225 85.340 ;
        RECT 136.575 85.140 152.225 85.340 ;
        RECT 152.575 85.140 154.225 85.340 ;
        RECT 6.890 84.740 7.290 85.140 ;
        RECT 8.890 84.740 9.290 85.140 ;
        RECT 10.890 84.740 11.290 85.140 ;
        RECT 12.890 84.740 13.290 85.140 ;
        RECT 14.890 84.740 15.290 85.140 ;
        RECT 16.890 84.740 17.290 85.140 ;
        RECT 18.890 84.740 19.290 85.140 ;
        RECT 20.890 84.740 21.290 85.140 ;
        RECT 22.890 84.740 23.290 85.140 ;
        RECT 24.890 84.740 25.290 85.140 ;
        RECT 26.890 84.740 27.290 85.140 ;
        RECT 28.890 84.740 29.290 85.140 ;
        RECT 30.890 84.740 31.290 85.140 ;
        RECT 32.890 84.740 33.290 85.140 ;
        RECT 34.890 84.740 35.290 85.140 ;
        RECT 36.890 84.740 37.290 85.140 ;
        RECT 38.890 84.740 39.290 85.140 ;
        RECT 40.890 84.740 41.290 85.140 ;
        RECT 42.890 84.740 43.290 85.140 ;
        RECT 44.890 84.740 45.290 85.140 ;
        RECT 46.890 84.740 47.290 85.140 ;
        RECT 48.890 84.740 49.290 85.140 ;
        RECT 50.890 84.740 51.290 85.140 ;
        RECT 52.890 84.740 53.290 85.140 ;
        RECT 54.890 84.740 55.290 85.140 ;
        RECT 56.890 84.740 57.290 85.140 ;
        RECT 58.890 84.740 59.290 85.140 ;
        RECT 60.890 84.740 61.290 85.140 ;
        RECT 62.890 84.740 63.290 85.140 ;
        RECT 64.890 84.740 65.290 85.140 ;
        RECT 66.890 84.740 67.290 85.140 ;
        RECT 68.890 84.740 69.290 85.140 ;
        RECT 70.890 84.740 71.290 85.140 ;
        RECT 72.890 84.740 73.290 85.140 ;
        RECT 87.825 84.740 88.225 85.140 ;
        RECT 89.825 84.740 90.225 85.140 ;
        RECT 91.825 84.740 92.225 85.140 ;
        RECT 93.825 84.740 94.225 85.140 ;
        RECT 95.825 84.740 96.225 85.140 ;
        RECT 97.825 84.740 98.225 85.140 ;
        RECT 99.825 84.740 100.225 85.140 ;
        RECT 101.825 84.740 102.225 85.140 ;
        RECT 103.825 84.740 104.225 85.140 ;
        RECT 105.825 84.740 106.225 85.140 ;
        RECT 107.825 84.740 108.225 85.140 ;
        RECT 109.825 84.740 110.225 85.140 ;
        RECT 111.825 84.740 112.225 85.140 ;
        RECT 113.825 84.740 114.225 85.140 ;
        RECT 115.825 84.740 116.225 85.140 ;
        RECT 117.825 84.740 118.225 85.140 ;
        RECT 119.825 84.740 120.225 85.140 ;
        RECT 121.825 84.740 122.225 85.140 ;
        RECT 123.825 84.740 124.225 85.140 ;
        RECT 125.825 84.740 126.225 85.140 ;
        RECT 127.825 84.740 128.225 85.140 ;
        RECT 129.825 84.740 130.225 85.140 ;
        RECT 131.825 84.740 132.225 85.140 ;
        RECT 133.825 84.740 134.225 85.140 ;
        RECT 135.825 84.740 136.225 85.140 ;
        RECT 137.825 84.740 138.225 85.140 ;
        RECT 139.825 84.740 140.225 85.140 ;
        RECT 141.825 84.740 142.225 85.140 ;
        RECT 143.825 84.740 144.225 85.140 ;
        RECT 145.825 84.740 146.225 85.140 ;
        RECT 147.825 84.740 148.225 85.140 ;
        RECT 149.825 84.740 150.225 85.140 ;
        RECT 151.825 84.740 152.225 85.140 ;
        RECT 153.825 84.740 154.225 85.140 ;
        RECT 6.960 83.890 7.220 84.740 ;
        RECT 8.990 83.890 9.190 84.740 ;
        RECT 10.990 83.890 11.190 84.740 ;
        RECT 12.990 83.890 13.190 84.740 ;
        RECT 14.990 83.890 15.190 84.740 ;
        RECT 16.990 83.890 17.190 84.740 ;
        RECT 18.990 83.890 19.190 84.740 ;
        RECT 20.990 83.890 21.190 84.740 ;
        RECT 22.990 83.890 23.190 84.740 ;
        RECT 24.990 83.890 25.190 84.740 ;
        RECT 26.990 83.890 27.190 84.740 ;
        RECT 28.990 83.890 29.190 84.740 ;
        RECT 30.990 83.890 31.190 84.740 ;
        RECT 32.990 83.890 33.190 84.740 ;
        RECT 34.990 83.890 35.190 84.740 ;
        RECT 36.990 83.890 37.190 84.740 ;
        RECT 38.990 83.890 39.190 84.740 ;
        RECT 40.990 83.890 41.190 84.740 ;
        RECT 42.990 83.890 43.190 84.740 ;
        RECT 44.990 83.890 45.190 84.740 ;
        RECT 46.990 83.890 47.190 84.740 ;
        RECT 113.925 83.890 114.125 84.740 ;
        RECT 115.925 83.890 116.125 84.740 ;
        RECT 117.925 83.890 118.125 84.740 ;
        RECT 119.925 83.890 120.125 84.740 ;
        RECT 121.925 83.890 122.125 84.740 ;
        RECT 123.925 83.890 124.125 84.740 ;
        RECT 125.925 83.890 126.125 84.740 ;
        RECT 127.925 83.890 128.125 84.740 ;
        RECT 129.925 83.890 130.125 84.740 ;
        RECT 131.925 83.890 132.125 84.740 ;
        RECT 133.925 83.890 134.125 84.740 ;
        RECT 135.925 83.890 136.125 84.740 ;
        RECT 137.925 83.890 138.125 84.740 ;
        RECT 139.925 83.890 140.125 84.740 ;
        RECT 141.925 83.890 142.125 84.740 ;
        RECT 143.925 83.890 144.125 84.740 ;
        RECT 145.925 83.890 146.125 84.740 ;
        RECT 147.925 83.890 148.125 84.740 ;
        RECT 149.925 83.890 150.125 84.740 ;
        RECT 151.925 83.890 152.125 84.740 ;
        RECT 153.895 83.890 154.155 84.740 ;
        RECT 6.890 83.490 7.290 83.890 ;
        RECT 8.890 83.490 9.290 83.890 ;
        RECT 10.890 83.490 11.290 83.890 ;
        RECT 12.890 83.490 13.290 83.890 ;
        RECT 14.890 83.490 15.290 83.890 ;
        RECT 16.890 83.490 17.290 83.890 ;
        RECT 18.890 83.490 19.290 83.890 ;
        RECT 20.890 83.490 21.290 83.890 ;
        RECT 22.890 83.490 23.290 83.890 ;
        RECT 24.890 83.490 25.290 83.890 ;
        RECT 26.890 83.490 27.290 83.890 ;
        RECT 28.890 83.490 29.290 83.890 ;
        RECT 30.890 83.490 31.290 83.890 ;
        RECT 32.890 83.490 33.290 83.890 ;
        RECT 34.890 83.490 35.290 83.890 ;
        RECT 36.890 83.490 37.290 83.890 ;
        RECT 38.890 83.490 39.290 83.890 ;
        RECT 40.890 83.490 41.290 83.890 ;
        RECT 42.890 83.490 43.290 83.890 ;
        RECT 44.890 83.490 45.290 83.890 ;
        RECT 46.890 83.490 47.290 83.890 ;
        RECT 48.890 83.490 49.290 83.890 ;
        RECT 50.890 83.490 51.290 83.890 ;
        RECT 52.890 83.490 53.290 83.890 ;
        RECT 54.890 83.490 55.290 83.890 ;
        RECT 56.890 83.490 57.290 83.890 ;
        RECT 58.890 83.490 59.290 83.890 ;
        RECT 60.890 83.490 61.290 83.890 ;
        RECT 62.890 83.490 63.290 83.890 ;
        RECT 64.890 83.490 65.290 83.890 ;
        RECT 66.890 83.490 67.290 83.890 ;
        RECT 68.890 83.490 69.290 83.890 ;
        RECT 70.890 83.490 71.290 83.890 ;
        RECT 72.890 83.490 73.290 83.890 ;
        RECT 87.825 83.490 88.225 83.890 ;
        RECT 89.825 83.490 90.225 83.890 ;
        RECT 91.825 83.490 92.225 83.890 ;
        RECT 93.825 83.490 94.225 83.890 ;
        RECT 95.825 83.490 96.225 83.890 ;
        RECT 97.825 83.490 98.225 83.890 ;
        RECT 99.825 83.490 100.225 83.890 ;
        RECT 101.825 83.490 102.225 83.890 ;
        RECT 103.825 83.490 104.225 83.890 ;
        RECT 105.825 83.490 106.225 83.890 ;
        RECT 107.825 83.490 108.225 83.890 ;
        RECT 109.825 83.490 110.225 83.890 ;
        RECT 111.825 83.490 112.225 83.890 ;
        RECT 113.825 83.490 114.225 83.890 ;
        RECT 115.825 83.490 116.225 83.890 ;
        RECT 117.825 83.490 118.225 83.890 ;
        RECT 119.825 83.490 120.225 83.890 ;
        RECT 121.825 83.490 122.225 83.890 ;
        RECT 123.825 83.490 124.225 83.890 ;
        RECT 125.825 83.490 126.225 83.890 ;
        RECT 127.825 83.490 128.225 83.890 ;
        RECT 129.825 83.490 130.225 83.890 ;
        RECT 131.825 83.490 132.225 83.890 ;
        RECT 133.825 83.490 134.225 83.890 ;
        RECT 135.825 83.490 136.225 83.890 ;
        RECT 137.825 83.490 138.225 83.890 ;
        RECT 139.825 83.490 140.225 83.890 ;
        RECT 141.825 83.490 142.225 83.890 ;
        RECT 143.825 83.490 144.225 83.890 ;
        RECT 145.825 83.490 146.225 83.890 ;
        RECT 147.825 83.490 148.225 83.890 ;
        RECT 149.825 83.490 150.225 83.890 ;
        RECT 151.825 83.490 152.225 83.890 ;
        RECT 153.825 83.490 154.225 83.890 ;
        RECT 6.890 83.290 8.540 83.490 ;
        RECT 8.890 83.290 24.540 83.490 ;
        RECT 24.890 83.290 38.540 83.490 ;
        RECT 38.890 83.290 48.540 83.490 ;
        RECT 48.890 83.290 74.540 83.490 ;
        RECT 86.575 83.290 112.225 83.490 ;
        RECT 112.575 83.290 122.225 83.490 ;
        RECT 122.575 83.290 136.225 83.490 ;
        RECT 136.575 83.290 152.225 83.490 ;
        RECT 152.575 83.290 154.225 83.490 ;
        RECT 6.890 82.890 7.290 83.290 ;
        RECT 8.890 82.890 9.290 83.290 ;
        RECT 10.890 82.890 11.290 83.290 ;
        RECT 12.890 82.890 13.290 83.290 ;
        RECT 14.890 82.890 15.290 83.290 ;
        RECT 16.890 82.890 17.290 83.290 ;
        RECT 18.890 82.890 19.290 83.290 ;
        RECT 20.890 82.890 21.290 83.290 ;
        RECT 22.890 82.890 23.290 83.290 ;
        RECT 24.890 82.890 25.290 83.290 ;
        RECT 26.890 82.890 27.290 83.290 ;
        RECT 28.890 82.890 29.290 83.290 ;
        RECT 30.890 82.890 31.290 83.290 ;
        RECT 32.890 82.890 33.290 83.290 ;
        RECT 34.890 82.890 35.290 83.290 ;
        RECT 36.890 82.890 37.290 83.290 ;
        RECT 38.890 82.890 39.290 83.290 ;
        RECT 40.890 82.890 41.290 83.290 ;
        RECT 42.890 82.890 43.290 83.290 ;
        RECT 44.890 82.890 45.290 83.290 ;
        RECT 46.890 82.890 47.290 83.290 ;
        RECT 48.890 82.890 49.290 83.290 ;
        RECT 50.890 82.890 51.290 83.290 ;
        RECT 52.890 82.890 53.290 83.290 ;
        RECT 54.890 82.890 55.290 83.290 ;
        RECT 56.890 82.890 57.290 83.290 ;
        RECT 58.890 82.890 59.290 83.290 ;
        RECT 60.890 82.890 61.290 83.290 ;
        RECT 62.890 82.890 63.290 83.290 ;
        RECT 64.890 82.890 65.290 83.290 ;
        RECT 66.890 82.890 67.290 83.290 ;
        RECT 68.890 82.890 69.290 83.290 ;
        RECT 70.890 82.890 71.290 83.290 ;
        RECT 72.890 82.890 73.290 83.290 ;
        RECT 87.825 82.890 88.225 83.290 ;
        RECT 89.825 82.890 90.225 83.290 ;
        RECT 91.825 82.890 92.225 83.290 ;
        RECT 93.825 82.890 94.225 83.290 ;
        RECT 95.825 82.890 96.225 83.290 ;
        RECT 97.825 82.890 98.225 83.290 ;
        RECT 99.825 82.890 100.225 83.290 ;
        RECT 101.825 82.890 102.225 83.290 ;
        RECT 103.825 82.890 104.225 83.290 ;
        RECT 105.825 82.890 106.225 83.290 ;
        RECT 107.825 82.890 108.225 83.290 ;
        RECT 109.825 82.890 110.225 83.290 ;
        RECT 111.825 82.890 112.225 83.290 ;
        RECT 113.825 82.890 114.225 83.290 ;
        RECT 115.825 82.890 116.225 83.290 ;
        RECT 117.825 82.890 118.225 83.290 ;
        RECT 119.825 82.890 120.225 83.290 ;
        RECT 121.825 82.890 122.225 83.290 ;
        RECT 123.825 82.890 124.225 83.290 ;
        RECT 125.825 82.890 126.225 83.290 ;
        RECT 127.825 82.890 128.225 83.290 ;
        RECT 129.825 82.890 130.225 83.290 ;
        RECT 131.825 82.890 132.225 83.290 ;
        RECT 133.825 82.890 134.225 83.290 ;
        RECT 135.825 82.890 136.225 83.290 ;
        RECT 137.825 82.890 138.225 83.290 ;
        RECT 139.825 82.890 140.225 83.290 ;
        RECT 141.825 82.890 142.225 83.290 ;
        RECT 143.825 82.890 144.225 83.290 ;
        RECT 145.825 82.890 146.225 83.290 ;
        RECT 147.825 82.890 148.225 83.290 ;
        RECT 149.825 82.890 150.225 83.290 ;
        RECT 151.825 82.890 152.225 83.290 ;
        RECT 153.825 82.890 154.225 83.290 ;
        RECT 6.960 82.040 7.220 82.890 ;
        RECT 8.990 82.040 9.190 82.890 ;
        RECT 10.990 82.040 11.190 82.890 ;
        RECT 12.990 82.040 13.190 82.890 ;
        RECT 14.990 82.040 15.190 82.890 ;
        RECT 16.990 82.040 17.190 82.890 ;
        RECT 18.990 82.040 19.190 82.890 ;
        RECT 20.990 82.040 21.190 82.890 ;
        RECT 22.990 82.040 23.190 82.890 ;
        RECT 24.990 82.040 25.190 82.890 ;
        RECT 26.990 82.040 27.190 82.890 ;
        RECT 28.990 82.040 29.190 82.890 ;
        RECT 30.990 82.040 31.190 82.890 ;
        RECT 32.990 82.040 33.190 82.890 ;
        RECT 34.990 82.040 35.190 82.890 ;
        RECT 36.990 82.040 37.190 82.890 ;
        RECT 38.990 82.040 39.190 82.890 ;
        RECT 40.990 82.040 41.190 82.890 ;
        RECT 42.990 82.040 43.190 82.890 ;
        RECT 44.990 82.040 45.190 82.890 ;
        RECT 46.990 82.040 47.190 82.890 ;
        RECT 48.990 82.040 49.190 82.890 ;
        RECT 50.990 82.040 51.190 82.890 ;
        RECT 52.990 82.040 53.190 82.890 ;
        RECT 54.990 82.040 55.190 82.890 ;
        RECT 56.990 82.040 57.190 82.890 ;
        RECT 58.990 82.040 59.190 82.890 ;
        RECT 60.990 82.040 61.190 82.890 ;
        RECT 62.990 82.040 63.190 82.890 ;
        RECT 64.990 82.040 65.190 82.890 ;
        RECT 66.990 82.040 67.190 82.890 ;
        RECT 68.990 82.040 69.190 82.890 ;
        RECT 70.990 82.040 71.190 82.890 ;
        RECT 89.925 82.040 90.125 82.890 ;
        RECT 91.925 82.040 92.125 82.890 ;
        RECT 93.925 82.040 94.125 82.890 ;
        RECT 95.925 82.040 96.125 82.890 ;
        RECT 97.925 82.040 98.125 82.890 ;
        RECT 99.925 82.040 100.125 82.890 ;
        RECT 101.925 82.040 102.125 82.890 ;
        RECT 103.925 82.040 104.125 82.890 ;
        RECT 105.925 82.040 106.125 82.890 ;
        RECT 107.925 82.040 108.125 82.890 ;
        RECT 109.925 82.040 110.125 82.890 ;
        RECT 111.925 82.040 112.125 82.890 ;
        RECT 113.925 82.040 114.125 82.890 ;
        RECT 115.925 82.040 116.125 82.890 ;
        RECT 117.925 82.040 118.125 82.890 ;
        RECT 119.925 82.040 120.125 82.890 ;
        RECT 121.925 82.040 122.125 82.890 ;
        RECT 123.925 82.040 124.125 82.890 ;
        RECT 125.925 82.040 126.125 82.890 ;
        RECT 127.925 82.040 128.125 82.890 ;
        RECT 129.925 82.040 130.125 82.890 ;
        RECT 131.925 82.040 132.125 82.890 ;
        RECT 133.925 82.040 134.125 82.890 ;
        RECT 135.925 82.040 136.125 82.890 ;
        RECT 137.925 82.040 138.125 82.890 ;
        RECT 139.925 82.040 140.125 82.890 ;
        RECT 141.925 82.040 142.125 82.890 ;
        RECT 143.925 82.040 144.125 82.890 ;
        RECT 145.925 82.040 146.125 82.890 ;
        RECT 147.925 82.040 148.125 82.890 ;
        RECT 149.925 82.040 150.125 82.890 ;
        RECT 151.925 82.040 152.125 82.890 ;
        RECT 153.895 82.040 154.155 82.890 ;
        RECT 6.890 81.640 7.290 82.040 ;
        RECT 8.890 81.640 9.290 82.040 ;
        RECT 10.890 81.640 11.290 82.040 ;
        RECT 12.890 81.640 13.290 82.040 ;
        RECT 14.890 81.640 15.290 82.040 ;
        RECT 16.890 81.640 17.290 82.040 ;
        RECT 18.890 81.640 19.290 82.040 ;
        RECT 20.890 81.640 21.290 82.040 ;
        RECT 22.890 81.640 23.290 82.040 ;
        RECT 24.890 81.640 25.290 82.040 ;
        RECT 26.890 81.640 27.290 82.040 ;
        RECT 28.890 81.640 29.290 82.040 ;
        RECT 30.890 81.640 31.290 82.040 ;
        RECT 32.890 81.640 33.290 82.040 ;
        RECT 34.890 81.640 35.290 82.040 ;
        RECT 36.890 81.640 37.290 82.040 ;
        RECT 38.890 81.640 39.290 82.040 ;
        RECT 40.890 81.640 41.290 82.040 ;
        RECT 42.890 81.640 43.290 82.040 ;
        RECT 44.890 81.640 45.290 82.040 ;
        RECT 46.890 81.640 47.290 82.040 ;
        RECT 48.890 81.640 49.290 82.040 ;
        RECT 50.890 81.640 51.290 82.040 ;
        RECT 52.890 81.640 53.290 82.040 ;
        RECT 54.890 81.640 55.290 82.040 ;
        RECT 56.890 81.640 57.290 82.040 ;
        RECT 58.890 81.640 59.290 82.040 ;
        RECT 60.890 81.640 61.290 82.040 ;
        RECT 62.890 81.640 63.290 82.040 ;
        RECT 64.890 81.640 65.290 82.040 ;
        RECT 66.890 81.640 67.290 82.040 ;
        RECT 68.890 81.640 69.290 82.040 ;
        RECT 70.890 81.640 71.290 82.040 ;
        RECT 72.890 81.640 73.290 82.040 ;
        RECT 87.825 81.640 88.225 82.040 ;
        RECT 89.825 81.640 90.225 82.040 ;
        RECT 91.825 81.640 92.225 82.040 ;
        RECT 93.825 81.640 94.225 82.040 ;
        RECT 95.825 81.640 96.225 82.040 ;
        RECT 97.825 81.640 98.225 82.040 ;
        RECT 99.825 81.640 100.225 82.040 ;
        RECT 101.825 81.640 102.225 82.040 ;
        RECT 103.825 81.640 104.225 82.040 ;
        RECT 105.825 81.640 106.225 82.040 ;
        RECT 107.825 81.640 108.225 82.040 ;
        RECT 109.825 81.640 110.225 82.040 ;
        RECT 111.825 81.640 112.225 82.040 ;
        RECT 113.825 81.640 114.225 82.040 ;
        RECT 115.825 81.640 116.225 82.040 ;
        RECT 117.825 81.640 118.225 82.040 ;
        RECT 119.825 81.640 120.225 82.040 ;
        RECT 121.825 81.640 122.225 82.040 ;
        RECT 123.825 81.640 124.225 82.040 ;
        RECT 125.825 81.640 126.225 82.040 ;
        RECT 127.825 81.640 128.225 82.040 ;
        RECT 129.825 81.640 130.225 82.040 ;
        RECT 131.825 81.640 132.225 82.040 ;
        RECT 133.825 81.640 134.225 82.040 ;
        RECT 135.825 81.640 136.225 82.040 ;
        RECT 137.825 81.640 138.225 82.040 ;
        RECT 139.825 81.640 140.225 82.040 ;
        RECT 141.825 81.640 142.225 82.040 ;
        RECT 143.825 81.640 144.225 82.040 ;
        RECT 145.825 81.640 146.225 82.040 ;
        RECT 147.825 81.640 148.225 82.040 ;
        RECT 149.825 81.640 150.225 82.040 ;
        RECT 151.825 81.640 152.225 82.040 ;
        RECT 153.825 81.640 154.225 82.040 ;
        RECT 6.890 81.440 8.540 81.640 ;
        RECT 8.890 81.440 24.540 81.640 ;
        RECT 24.890 81.440 38.540 81.640 ;
        RECT 38.890 81.440 48.540 81.640 ;
        RECT 48.890 81.440 74.540 81.640 ;
        RECT 86.575 81.440 112.225 81.640 ;
        RECT 112.575 81.440 122.225 81.640 ;
        RECT 122.575 81.440 136.225 81.640 ;
        RECT 136.575 81.440 152.225 81.640 ;
        RECT 152.575 81.440 154.225 81.640 ;
        RECT 6.890 81.040 7.290 81.440 ;
        RECT 8.890 81.040 9.290 81.440 ;
        RECT 10.890 81.040 11.290 81.440 ;
        RECT 12.890 81.040 13.290 81.440 ;
        RECT 14.890 81.040 15.290 81.440 ;
        RECT 16.890 81.040 17.290 81.440 ;
        RECT 18.890 81.040 19.290 81.440 ;
        RECT 20.890 81.040 21.290 81.440 ;
        RECT 22.890 81.040 23.290 81.440 ;
        RECT 24.890 81.040 25.290 81.440 ;
        RECT 26.890 81.040 27.290 81.440 ;
        RECT 28.890 81.040 29.290 81.440 ;
        RECT 30.890 81.040 31.290 81.440 ;
        RECT 32.890 81.040 33.290 81.440 ;
        RECT 34.890 81.040 35.290 81.440 ;
        RECT 36.890 81.040 37.290 81.440 ;
        RECT 38.890 81.040 39.290 81.440 ;
        RECT 40.890 81.040 41.290 81.440 ;
        RECT 42.890 81.040 43.290 81.440 ;
        RECT 44.890 81.040 45.290 81.440 ;
        RECT 46.890 81.040 47.290 81.440 ;
        RECT 48.890 81.040 49.290 81.440 ;
        RECT 50.890 81.040 51.290 81.440 ;
        RECT 52.890 81.040 53.290 81.440 ;
        RECT 54.890 81.040 55.290 81.440 ;
        RECT 56.890 81.040 57.290 81.440 ;
        RECT 58.890 81.040 59.290 81.440 ;
        RECT 60.890 81.040 61.290 81.440 ;
        RECT 62.890 81.040 63.290 81.440 ;
        RECT 64.890 81.040 65.290 81.440 ;
        RECT 66.890 81.040 67.290 81.440 ;
        RECT 68.890 81.040 69.290 81.440 ;
        RECT 70.890 81.040 71.290 81.440 ;
        RECT 72.890 81.040 73.290 81.440 ;
        RECT 87.825 81.040 88.225 81.440 ;
        RECT 89.825 81.040 90.225 81.440 ;
        RECT 91.825 81.040 92.225 81.440 ;
        RECT 93.825 81.040 94.225 81.440 ;
        RECT 95.825 81.040 96.225 81.440 ;
        RECT 97.825 81.040 98.225 81.440 ;
        RECT 99.825 81.040 100.225 81.440 ;
        RECT 101.825 81.040 102.225 81.440 ;
        RECT 103.825 81.040 104.225 81.440 ;
        RECT 105.825 81.040 106.225 81.440 ;
        RECT 107.825 81.040 108.225 81.440 ;
        RECT 109.825 81.040 110.225 81.440 ;
        RECT 111.825 81.040 112.225 81.440 ;
        RECT 113.825 81.040 114.225 81.440 ;
        RECT 115.825 81.040 116.225 81.440 ;
        RECT 117.825 81.040 118.225 81.440 ;
        RECT 119.825 81.040 120.225 81.440 ;
        RECT 121.825 81.040 122.225 81.440 ;
        RECT 123.825 81.040 124.225 81.440 ;
        RECT 125.825 81.040 126.225 81.440 ;
        RECT 127.825 81.040 128.225 81.440 ;
        RECT 129.825 81.040 130.225 81.440 ;
        RECT 131.825 81.040 132.225 81.440 ;
        RECT 133.825 81.040 134.225 81.440 ;
        RECT 135.825 81.040 136.225 81.440 ;
        RECT 137.825 81.040 138.225 81.440 ;
        RECT 139.825 81.040 140.225 81.440 ;
        RECT 141.825 81.040 142.225 81.440 ;
        RECT 143.825 81.040 144.225 81.440 ;
        RECT 145.825 81.040 146.225 81.440 ;
        RECT 147.825 81.040 148.225 81.440 ;
        RECT 149.825 81.040 150.225 81.440 ;
        RECT 151.825 81.040 152.225 81.440 ;
        RECT 153.825 81.040 154.225 81.440 ;
        RECT 6.960 80.190 7.220 81.040 ;
        RECT 8.990 80.190 9.190 81.040 ;
        RECT 10.990 80.190 11.190 81.040 ;
        RECT 12.990 80.190 13.190 81.040 ;
        RECT 14.990 80.190 15.190 81.040 ;
        RECT 16.990 80.190 17.190 81.040 ;
        RECT 18.990 80.190 19.190 81.040 ;
        RECT 20.990 80.190 21.190 81.040 ;
        RECT 24.990 80.190 25.190 81.040 ;
        RECT 26.990 80.190 27.190 81.040 ;
        RECT 28.990 80.190 29.190 81.040 ;
        RECT 30.990 80.190 31.190 81.040 ;
        RECT 32.990 80.190 33.190 81.040 ;
        RECT 34.990 80.190 35.190 81.040 ;
        RECT 36.990 80.190 37.190 81.040 ;
        RECT 38.990 80.190 39.190 81.040 ;
        RECT 40.990 80.190 41.190 81.040 ;
        RECT 42.990 80.190 43.190 81.040 ;
        RECT 44.990 80.190 45.190 81.040 ;
        RECT 48.990 80.190 49.190 81.040 ;
        RECT 50.990 80.190 51.190 81.040 ;
        RECT 52.990 80.190 53.190 81.040 ;
        RECT 54.990 80.190 55.190 81.040 ;
        RECT 56.990 80.190 57.190 81.040 ;
        RECT 58.990 80.190 59.190 81.040 ;
        RECT 60.990 80.190 61.190 81.040 ;
        RECT 62.990 80.190 63.190 81.040 ;
        RECT 64.990 80.190 65.190 81.040 ;
        RECT 66.990 80.190 67.190 81.040 ;
        RECT 68.990 80.190 69.190 81.040 ;
        RECT 70.990 80.190 71.190 81.040 ;
        RECT 89.925 80.190 90.125 81.040 ;
        RECT 91.925 80.190 92.125 81.040 ;
        RECT 93.925 80.190 94.125 81.040 ;
        RECT 95.925 80.190 96.125 81.040 ;
        RECT 97.925 80.190 98.125 81.040 ;
        RECT 99.925 80.190 100.125 81.040 ;
        RECT 101.925 80.190 102.125 81.040 ;
        RECT 103.925 80.190 104.125 81.040 ;
        RECT 105.925 80.190 106.125 81.040 ;
        RECT 107.925 80.190 108.125 81.040 ;
        RECT 109.925 80.190 110.125 81.040 ;
        RECT 111.925 80.190 112.125 81.040 ;
        RECT 115.925 80.190 116.125 81.040 ;
        RECT 117.925 80.190 118.125 81.040 ;
        RECT 119.925 80.190 120.125 81.040 ;
        RECT 121.925 80.190 122.125 81.040 ;
        RECT 123.925 80.190 124.125 81.040 ;
        RECT 125.925 80.190 126.125 81.040 ;
        RECT 127.925 80.190 128.125 81.040 ;
        RECT 129.925 80.190 130.125 81.040 ;
        RECT 131.925 80.190 132.125 81.040 ;
        RECT 133.925 80.190 134.125 81.040 ;
        RECT 135.925 80.190 136.125 81.040 ;
        RECT 139.925 80.190 140.125 81.040 ;
        RECT 141.925 80.190 142.125 81.040 ;
        RECT 143.925 80.190 144.125 81.040 ;
        RECT 145.925 80.190 146.125 81.040 ;
        RECT 147.925 80.190 148.125 81.040 ;
        RECT 149.925 80.190 150.125 81.040 ;
        RECT 151.925 80.190 152.125 81.040 ;
        RECT 153.895 80.190 154.155 81.040 ;
        RECT 6.890 79.790 7.290 80.190 ;
        RECT 8.890 79.790 9.290 80.190 ;
        RECT 10.890 79.790 11.290 80.190 ;
        RECT 12.890 79.790 13.290 80.190 ;
        RECT 14.890 79.790 15.290 80.190 ;
        RECT 16.890 79.790 17.290 80.190 ;
        RECT 18.890 79.790 19.290 80.190 ;
        RECT 20.890 79.790 21.290 80.190 ;
        RECT 22.890 79.790 23.290 80.190 ;
        RECT 24.890 79.790 25.290 80.190 ;
        RECT 26.890 79.790 27.290 80.190 ;
        RECT 28.890 79.790 29.290 80.190 ;
        RECT 30.890 79.790 31.290 80.190 ;
        RECT 32.890 79.790 33.290 80.190 ;
        RECT 34.890 79.790 35.290 80.190 ;
        RECT 36.890 79.790 37.290 80.190 ;
        RECT 38.890 79.790 39.290 80.190 ;
        RECT 40.890 79.790 41.290 80.190 ;
        RECT 42.890 79.790 43.290 80.190 ;
        RECT 44.890 79.790 45.290 80.190 ;
        RECT 46.890 79.790 47.290 80.190 ;
        RECT 48.890 79.790 49.290 80.190 ;
        RECT 50.890 79.790 51.290 80.190 ;
        RECT 52.890 79.790 53.290 80.190 ;
        RECT 54.890 79.790 55.290 80.190 ;
        RECT 56.890 79.790 57.290 80.190 ;
        RECT 58.890 79.790 59.290 80.190 ;
        RECT 60.890 79.790 61.290 80.190 ;
        RECT 62.890 79.790 63.290 80.190 ;
        RECT 64.890 79.790 65.290 80.190 ;
        RECT 66.890 79.790 67.290 80.190 ;
        RECT 68.890 79.790 69.290 80.190 ;
        RECT 70.890 79.790 71.290 80.190 ;
        RECT 72.890 79.790 73.290 80.190 ;
        RECT 87.825 79.790 88.225 80.190 ;
        RECT 89.825 79.790 90.225 80.190 ;
        RECT 91.825 79.790 92.225 80.190 ;
        RECT 93.825 79.790 94.225 80.190 ;
        RECT 95.825 79.790 96.225 80.190 ;
        RECT 97.825 79.790 98.225 80.190 ;
        RECT 99.825 79.790 100.225 80.190 ;
        RECT 101.825 79.790 102.225 80.190 ;
        RECT 103.825 79.790 104.225 80.190 ;
        RECT 105.825 79.790 106.225 80.190 ;
        RECT 107.825 79.790 108.225 80.190 ;
        RECT 109.825 79.790 110.225 80.190 ;
        RECT 111.825 79.790 112.225 80.190 ;
        RECT 113.825 79.790 114.225 80.190 ;
        RECT 115.825 79.790 116.225 80.190 ;
        RECT 117.825 79.790 118.225 80.190 ;
        RECT 119.825 79.790 120.225 80.190 ;
        RECT 121.825 79.790 122.225 80.190 ;
        RECT 123.825 79.790 124.225 80.190 ;
        RECT 125.825 79.790 126.225 80.190 ;
        RECT 127.825 79.790 128.225 80.190 ;
        RECT 129.825 79.790 130.225 80.190 ;
        RECT 131.825 79.790 132.225 80.190 ;
        RECT 133.825 79.790 134.225 80.190 ;
        RECT 135.825 79.790 136.225 80.190 ;
        RECT 137.825 79.790 138.225 80.190 ;
        RECT 139.825 79.790 140.225 80.190 ;
        RECT 141.825 79.790 142.225 80.190 ;
        RECT 143.825 79.790 144.225 80.190 ;
        RECT 145.825 79.790 146.225 80.190 ;
        RECT 147.825 79.790 148.225 80.190 ;
        RECT 149.825 79.790 150.225 80.190 ;
        RECT 151.825 79.790 152.225 80.190 ;
        RECT 153.825 79.790 154.225 80.190 ;
        RECT 6.890 79.590 8.540 79.790 ;
        RECT 8.890 79.590 22.540 79.790 ;
        RECT 22.890 79.590 38.540 79.790 ;
        RECT 38.890 79.590 46.540 79.790 ;
        RECT 46.890 79.590 74.540 79.790 ;
        RECT 86.575 79.590 114.225 79.790 ;
        RECT 114.575 79.590 122.225 79.790 ;
        RECT 122.575 79.590 138.225 79.790 ;
        RECT 138.575 79.590 152.225 79.790 ;
        RECT 152.575 79.590 154.225 79.790 ;
        RECT 6.890 79.190 7.290 79.590 ;
        RECT 8.890 79.190 9.290 79.590 ;
        RECT 10.890 79.190 11.290 79.590 ;
        RECT 12.890 79.190 13.290 79.590 ;
        RECT 14.890 79.190 15.290 79.590 ;
        RECT 16.890 79.190 17.290 79.590 ;
        RECT 18.890 79.190 19.290 79.590 ;
        RECT 20.890 79.190 21.290 79.590 ;
        RECT 22.890 79.190 23.290 79.590 ;
        RECT 24.890 79.190 25.290 79.590 ;
        RECT 26.890 79.190 27.290 79.590 ;
        RECT 28.890 79.190 29.290 79.590 ;
        RECT 30.890 79.190 31.290 79.590 ;
        RECT 32.890 79.190 33.290 79.590 ;
        RECT 34.890 79.190 35.290 79.590 ;
        RECT 36.890 79.190 37.290 79.590 ;
        RECT 38.890 79.190 39.290 79.590 ;
        RECT 40.890 79.190 41.290 79.590 ;
        RECT 42.890 79.190 43.290 79.590 ;
        RECT 44.890 79.190 45.290 79.590 ;
        RECT 46.890 79.190 47.290 79.590 ;
        RECT 48.890 79.190 49.290 79.590 ;
        RECT 50.890 79.190 51.290 79.590 ;
        RECT 52.890 79.190 53.290 79.590 ;
        RECT 54.890 79.190 55.290 79.590 ;
        RECT 56.890 79.190 57.290 79.590 ;
        RECT 58.890 79.190 59.290 79.590 ;
        RECT 60.890 79.190 61.290 79.590 ;
        RECT 62.890 79.190 63.290 79.590 ;
        RECT 64.890 79.190 65.290 79.590 ;
        RECT 66.890 79.190 67.290 79.590 ;
        RECT 68.890 79.190 69.290 79.590 ;
        RECT 70.890 79.190 71.290 79.590 ;
        RECT 72.890 79.190 73.290 79.590 ;
        RECT 87.825 79.190 88.225 79.590 ;
        RECT 89.825 79.190 90.225 79.590 ;
        RECT 91.825 79.190 92.225 79.590 ;
        RECT 93.825 79.190 94.225 79.590 ;
        RECT 95.825 79.190 96.225 79.590 ;
        RECT 97.825 79.190 98.225 79.590 ;
        RECT 99.825 79.190 100.225 79.590 ;
        RECT 101.825 79.190 102.225 79.590 ;
        RECT 103.825 79.190 104.225 79.590 ;
        RECT 105.825 79.190 106.225 79.590 ;
        RECT 107.825 79.190 108.225 79.590 ;
        RECT 109.825 79.190 110.225 79.590 ;
        RECT 111.825 79.190 112.225 79.590 ;
        RECT 113.825 79.190 114.225 79.590 ;
        RECT 115.825 79.190 116.225 79.590 ;
        RECT 117.825 79.190 118.225 79.590 ;
        RECT 119.825 79.190 120.225 79.590 ;
        RECT 121.825 79.190 122.225 79.590 ;
        RECT 123.825 79.190 124.225 79.590 ;
        RECT 125.825 79.190 126.225 79.590 ;
        RECT 127.825 79.190 128.225 79.590 ;
        RECT 129.825 79.190 130.225 79.590 ;
        RECT 131.825 79.190 132.225 79.590 ;
        RECT 133.825 79.190 134.225 79.590 ;
        RECT 135.825 79.190 136.225 79.590 ;
        RECT 137.825 79.190 138.225 79.590 ;
        RECT 139.825 79.190 140.225 79.590 ;
        RECT 141.825 79.190 142.225 79.590 ;
        RECT 143.825 79.190 144.225 79.590 ;
        RECT 145.825 79.190 146.225 79.590 ;
        RECT 147.825 79.190 148.225 79.590 ;
        RECT 149.825 79.190 150.225 79.590 ;
        RECT 151.825 79.190 152.225 79.590 ;
        RECT 153.825 79.190 154.225 79.590 ;
        RECT 6.960 78.340 7.220 79.190 ;
        RECT 8.990 78.340 9.190 79.190 ;
        RECT 10.990 78.340 11.190 79.190 ;
        RECT 12.990 78.340 13.190 79.190 ;
        RECT 14.990 78.340 15.190 79.190 ;
        RECT 16.990 78.340 17.190 79.190 ;
        RECT 18.990 78.340 19.190 79.190 ;
        RECT 20.990 78.340 21.190 79.190 ;
        RECT 22.990 78.340 23.190 79.190 ;
        RECT 24.990 78.340 25.190 79.190 ;
        RECT 26.990 78.340 27.190 79.190 ;
        RECT 28.990 78.340 29.190 79.190 ;
        RECT 30.990 78.340 31.190 79.190 ;
        RECT 32.990 78.340 33.190 79.190 ;
        RECT 34.990 78.340 35.190 79.190 ;
        RECT 36.990 78.340 37.190 79.190 ;
        RECT 38.990 78.340 39.190 79.190 ;
        RECT 40.990 78.340 41.190 79.190 ;
        RECT 42.990 78.340 43.190 79.190 ;
        RECT 44.990 78.340 45.190 79.190 ;
        RECT 46.990 78.340 47.190 79.190 ;
        RECT 48.990 78.340 49.190 79.190 ;
        RECT 50.990 78.340 51.190 79.190 ;
        RECT 52.990 78.340 53.190 79.190 ;
        RECT 107.925 78.340 108.125 79.190 ;
        RECT 109.925 78.340 110.125 79.190 ;
        RECT 111.925 78.340 112.125 79.190 ;
        RECT 113.925 78.340 114.125 79.190 ;
        RECT 115.925 78.340 116.125 79.190 ;
        RECT 117.925 78.340 118.125 79.190 ;
        RECT 119.925 78.340 120.125 79.190 ;
        RECT 121.925 78.340 122.125 79.190 ;
        RECT 123.925 78.340 124.125 79.190 ;
        RECT 125.925 78.340 126.125 79.190 ;
        RECT 127.925 78.340 128.125 79.190 ;
        RECT 129.925 78.340 130.125 79.190 ;
        RECT 131.925 78.340 132.125 79.190 ;
        RECT 133.925 78.340 134.125 79.190 ;
        RECT 135.925 78.340 136.125 79.190 ;
        RECT 137.925 78.340 138.125 79.190 ;
        RECT 139.925 78.340 140.125 79.190 ;
        RECT 141.925 78.340 142.125 79.190 ;
        RECT 143.925 78.340 144.125 79.190 ;
        RECT 145.925 78.340 146.125 79.190 ;
        RECT 147.925 78.340 148.125 79.190 ;
        RECT 149.925 78.340 150.125 79.190 ;
        RECT 151.925 78.340 152.125 79.190 ;
        RECT 153.895 78.340 154.155 79.190 ;
        RECT 6.890 77.940 7.290 78.340 ;
        RECT 8.890 77.940 9.290 78.340 ;
        RECT 10.890 77.940 11.290 78.340 ;
        RECT 12.890 77.940 13.290 78.340 ;
        RECT 14.890 77.940 15.290 78.340 ;
        RECT 16.890 77.940 17.290 78.340 ;
        RECT 18.890 77.940 19.290 78.340 ;
        RECT 20.890 77.940 21.290 78.340 ;
        RECT 22.890 77.940 23.290 78.340 ;
        RECT 24.890 77.940 25.290 78.340 ;
        RECT 26.890 77.940 27.290 78.340 ;
        RECT 28.890 77.940 29.290 78.340 ;
        RECT 30.890 77.940 31.290 78.340 ;
        RECT 32.890 77.940 33.290 78.340 ;
        RECT 34.890 77.940 35.290 78.340 ;
        RECT 36.890 77.940 37.290 78.340 ;
        RECT 38.890 77.940 39.290 78.340 ;
        RECT 40.890 77.940 41.290 78.340 ;
        RECT 42.890 77.940 43.290 78.340 ;
        RECT 44.890 77.940 45.290 78.340 ;
        RECT 46.890 77.940 47.290 78.340 ;
        RECT 48.890 77.940 49.290 78.340 ;
        RECT 50.890 77.940 51.290 78.340 ;
        RECT 52.890 77.940 53.290 78.340 ;
        RECT 54.890 77.940 55.290 78.340 ;
        RECT 56.890 77.940 57.290 78.340 ;
        RECT 58.890 77.940 59.290 78.340 ;
        RECT 60.890 77.940 61.290 78.340 ;
        RECT 62.890 77.940 63.290 78.340 ;
        RECT 64.890 77.940 65.290 78.340 ;
        RECT 66.890 77.940 67.290 78.340 ;
        RECT 68.890 77.940 69.290 78.340 ;
        RECT 70.890 77.940 71.290 78.340 ;
        RECT 72.890 77.940 73.290 78.340 ;
        RECT 87.825 77.940 88.225 78.340 ;
        RECT 89.825 77.940 90.225 78.340 ;
        RECT 91.825 77.940 92.225 78.340 ;
        RECT 93.825 77.940 94.225 78.340 ;
        RECT 95.825 77.940 96.225 78.340 ;
        RECT 97.825 77.940 98.225 78.340 ;
        RECT 99.825 77.940 100.225 78.340 ;
        RECT 101.825 77.940 102.225 78.340 ;
        RECT 103.825 77.940 104.225 78.340 ;
        RECT 105.825 77.940 106.225 78.340 ;
        RECT 107.825 77.940 108.225 78.340 ;
        RECT 109.825 77.940 110.225 78.340 ;
        RECT 111.825 77.940 112.225 78.340 ;
        RECT 113.825 77.940 114.225 78.340 ;
        RECT 115.825 77.940 116.225 78.340 ;
        RECT 117.825 77.940 118.225 78.340 ;
        RECT 119.825 77.940 120.225 78.340 ;
        RECT 121.825 77.940 122.225 78.340 ;
        RECT 123.825 77.940 124.225 78.340 ;
        RECT 125.825 77.940 126.225 78.340 ;
        RECT 127.825 77.940 128.225 78.340 ;
        RECT 129.825 77.940 130.225 78.340 ;
        RECT 131.825 77.940 132.225 78.340 ;
        RECT 133.825 77.940 134.225 78.340 ;
        RECT 135.825 77.940 136.225 78.340 ;
        RECT 137.825 77.940 138.225 78.340 ;
        RECT 139.825 77.940 140.225 78.340 ;
        RECT 141.825 77.940 142.225 78.340 ;
        RECT 143.825 77.940 144.225 78.340 ;
        RECT 145.825 77.940 146.225 78.340 ;
        RECT 147.825 77.940 148.225 78.340 ;
        RECT 149.825 77.940 150.225 78.340 ;
        RECT 151.825 77.940 152.225 78.340 ;
        RECT 153.825 77.940 154.225 78.340 ;
        RECT 6.890 77.740 8.540 77.940 ;
        RECT 8.890 77.740 22.540 77.940 ;
        RECT 22.890 77.740 38.540 77.940 ;
        RECT 38.890 77.740 46.540 77.940 ;
        RECT 46.890 77.740 50.540 77.940 ;
        RECT 50.890 77.740 52.540 77.940 ;
        RECT 52.890 77.740 54.540 77.940 ;
        RECT 54.890 77.740 74.540 77.940 ;
        RECT 86.575 77.740 106.225 77.940 ;
        RECT 106.575 77.740 108.225 77.940 ;
        RECT 108.575 77.740 110.225 77.940 ;
        RECT 110.575 77.740 114.225 77.940 ;
        RECT 114.575 77.740 122.225 77.940 ;
        RECT 122.575 77.740 138.225 77.940 ;
        RECT 138.575 77.740 152.225 77.940 ;
        RECT 152.575 77.740 154.225 77.940 ;
        RECT 6.890 77.340 7.290 77.740 ;
        RECT 8.890 77.340 9.290 77.740 ;
        RECT 10.890 77.340 11.290 77.740 ;
        RECT 12.890 77.340 13.290 77.740 ;
        RECT 14.890 77.340 15.290 77.740 ;
        RECT 16.890 77.340 17.290 77.740 ;
        RECT 18.890 77.340 19.290 77.740 ;
        RECT 20.890 77.340 21.290 77.740 ;
        RECT 22.890 77.340 23.290 77.740 ;
        RECT 24.890 77.340 25.290 77.740 ;
        RECT 26.890 77.340 27.290 77.740 ;
        RECT 28.890 77.340 29.290 77.740 ;
        RECT 30.890 77.340 31.290 77.740 ;
        RECT 32.890 77.340 33.290 77.740 ;
        RECT 34.890 77.340 35.290 77.740 ;
        RECT 36.890 77.340 37.290 77.740 ;
        RECT 38.890 77.340 39.290 77.740 ;
        RECT 40.890 77.340 41.290 77.740 ;
        RECT 42.890 77.340 43.290 77.740 ;
        RECT 44.890 77.340 45.290 77.740 ;
        RECT 46.890 77.340 47.290 77.740 ;
        RECT 48.890 77.340 49.290 77.740 ;
        RECT 50.890 77.340 51.290 77.740 ;
        RECT 52.890 77.340 53.290 77.740 ;
        RECT 54.890 77.340 55.290 77.740 ;
        RECT 56.890 77.340 57.290 77.740 ;
        RECT 58.890 77.340 59.290 77.740 ;
        RECT 60.890 77.340 61.290 77.740 ;
        RECT 62.890 77.340 63.290 77.740 ;
        RECT 64.890 77.340 65.290 77.740 ;
        RECT 66.890 77.340 67.290 77.740 ;
        RECT 68.890 77.340 69.290 77.740 ;
        RECT 70.890 77.340 71.290 77.740 ;
        RECT 72.890 77.340 73.290 77.740 ;
        RECT 87.825 77.340 88.225 77.740 ;
        RECT 89.825 77.340 90.225 77.740 ;
        RECT 91.825 77.340 92.225 77.740 ;
        RECT 93.825 77.340 94.225 77.740 ;
        RECT 95.825 77.340 96.225 77.740 ;
        RECT 97.825 77.340 98.225 77.740 ;
        RECT 99.825 77.340 100.225 77.740 ;
        RECT 101.825 77.340 102.225 77.740 ;
        RECT 103.825 77.340 104.225 77.740 ;
        RECT 105.825 77.340 106.225 77.740 ;
        RECT 107.825 77.340 108.225 77.740 ;
        RECT 109.825 77.340 110.225 77.740 ;
        RECT 111.825 77.340 112.225 77.740 ;
        RECT 113.825 77.340 114.225 77.740 ;
        RECT 115.825 77.340 116.225 77.740 ;
        RECT 117.825 77.340 118.225 77.740 ;
        RECT 119.825 77.340 120.225 77.740 ;
        RECT 121.825 77.340 122.225 77.740 ;
        RECT 123.825 77.340 124.225 77.740 ;
        RECT 125.825 77.340 126.225 77.740 ;
        RECT 127.825 77.340 128.225 77.740 ;
        RECT 129.825 77.340 130.225 77.740 ;
        RECT 131.825 77.340 132.225 77.740 ;
        RECT 133.825 77.340 134.225 77.740 ;
        RECT 135.825 77.340 136.225 77.740 ;
        RECT 137.825 77.340 138.225 77.740 ;
        RECT 139.825 77.340 140.225 77.740 ;
        RECT 141.825 77.340 142.225 77.740 ;
        RECT 143.825 77.340 144.225 77.740 ;
        RECT 145.825 77.340 146.225 77.740 ;
        RECT 147.825 77.340 148.225 77.740 ;
        RECT 149.825 77.340 150.225 77.740 ;
        RECT 151.825 77.340 152.225 77.740 ;
        RECT 153.825 77.340 154.225 77.740 ;
        RECT 6.960 76.490 7.220 77.340 ;
        RECT 8.990 76.490 9.190 77.340 ;
        RECT 10.990 76.490 11.190 77.340 ;
        RECT 12.990 76.490 13.190 77.340 ;
        RECT 14.990 76.490 15.190 77.340 ;
        RECT 16.990 76.490 17.190 77.340 ;
        RECT 18.990 76.490 19.190 77.340 ;
        RECT 20.990 76.490 21.190 77.340 ;
        RECT 22.990 76.490 23.190 77.340 ;
        RECT 24.990 76.490 25.190 77.340 ;
        RECT 26.990 76.490 27.190 77.340 ;
        RECT 28.990 76.490 29.190 77.340 ;
        RECT 30.990 76.490 31.190 77.340 ;
        RECT 32.990 76.490 33.190 77.340 ;
        RECT 34.990 76.490 35.190 77.340 ;
        RECT 36.990 76.490 37.190 77.340 ;
        RECT 38.990 76.490 39.190 77.340 ;
        RECT 40.990 76.490 41.190 77.340 ;
        RECT 42.990 76.490 43.190 77.340 ;
        RECT 44.990 76.490 45.190 77.340 ;
        RECT 46.990 76.490 47.190 77.340 ;
        RECT 48.990 76.490 49.190 77.340 ;
        RECT 50.990 76.490 51.190 77.340 ;
        RECT 52.990 76.490 53.190 77.340 ;
        RECT 54.990 76.490 55.190 77.340 ;
        RECT 56.990 76.490 57.190 77.340 ;
        RECT 58.990 76.490 59.190 77.340 ;
        RECT 60.990 76.490 61.190 77.340 ;
        RECT 62.990 76.490 63.190 77.340 ;
        RECT 64.990 76.490 65.190 77.340 ;
        RECT 66.990 76.490 67.190 77.340 ;
        RECT 68.990 76.490 69.190 77.340 ;
        RECT 70.990 76.490 71.190 77.340 ;
        RECT 89.925 76.490 90.125 77.340 ;
        RECT 91.925 76.490 92.125 77.340 ;
        RECT 93.925 76.490 94.125 77.340 ;
        RECT 95.925 76.490 96.125 77.340 ;
        RECT 97.925 76.490 98.125 77.340 ;
        RECT 99.925 76.490 100.125 77.340 ;
        RECT 101.925 76.490 102.125 77.340 ;
        RECT 103.925 76.490 104.125 77.340 ;
        RECT 105.925 76.490 106.125 77.340 ;
        RECT 107.925 76.490 108.125 77.340 ;
        RECT 109.925 76.490 110.125 77.340 ;
        RECT 111.925 76.490 112.125 77.340 ;
        RECT 113.925 76.490 114.125 77.340 ;
        RECT 115.925 76.490 116.125 77.340 ;
        RECT 117.925 76.490 118.125 77.340 ;
        RECT 119.925 76.490 120.125 77.340 ;
        RECT 121.925 76.490 122.125 77.340 ;
        RECT 123.925 76.490 124.125 77.340 ;
        RECT 125.925 76.490 126.125 77.340 ;
        RECT 127.925 76.490 128.125 77.340 ;
        RECT 129.925 76.490 130.125 77.340 ;
        RECT 131.925 76.490 132.125 77.340 ;
        RECT 133.925 76.490 134.125 77.340 ;
        RECT 135.925 76.490 136.125 77.340 ;
        RECT 137.925 76.490 138.125 77.340 ;
        RECT 139.925 76.490 140.125 77.340 ;
        RECT 141.925 76.490 142.125 77.340 ;
        RECT 143.925 76.490 144.125 77.340 ;
        RECT 145.925 76.490 146.125 77.340 ;
        RECT 147.925 76.490 148.125 77.340 ;
        RECT 149.925 76.490 150.125 77.340 ;
        RECT 151.925 76.490 152.125 77.340 ;
        RECT 153.895 76.490 154.155 77.340 ;
        RECT 6.890 76.090 7.290 76.490 ;
        RECT 8.890 76.090 9.290 76.490 ;
        RECT 10.890 76.090 11.290 76.490 ;
        RECT 12.890 76.090 13.290 76.490 ;
        RECT 14.890 76.090 15.290 76.490 ;
        RECT 16.890 76.090 17.290 76.490 ;
        RECT 18.890 76.090 19.290 76.490 ;
        RECT 20.890 76.090 21.290 76.490 ;
        RECT 22.890 76.090 23.290 76.490 ;
        RECT 24.890 76.090 25.290 76.490 ;
        RECT 26.890 76.090 27.290 76.490 ;
        RECT 28.890 76.090 29.290 76.490 ;
        RECT 30.890 76.090 31.290 76.490 ;
        RECT 32.890 76.090 33.290 76.490 ;
        RECT 34.890 76.090 35.290 76.490 ;
        RECT 36.890 76.090 37.290 76.490 ;
        RECT 38.890 76.090 39.290 76.490 ;
        RECT 40.890 76.090 41.290 76.490 ;
        RECT 42.890 76.090 43.290 76.490 ;
        RECT 44.890 76.090 45.290 76.490 ;
        RECT 46.890 76.090 47.290 76.490 ;
        RECT 48.890 76.090 49.290 76.490 ;
        RECT 50.890 76.090 51.290 76.490 ;
        RECT 52.890 76.090 53.290 76.490 ;
        RECT 54.890 76.090 55.290 76.490 ;
        RECT 56.890 76.090 57.290 76.490 ;
        RECT 58.890 76.090 59.290 76.490 ;
        RECT 60.890 76.090 61.290 76.490 ;
        RECT 62.890 76.090 63.290 76.490 ;
        RECT 64.890 76.090 65.290 76.490 ;
        RECT 66.890 76.090 67.290 76.490 ;
        RECT 68.890 76.090 69.290 76.490 ;
        RECT 70.890 76.090 71.290 76.490 ;
        RECT 72.890 76.090 73.290 76.490 ;
        RECT 87.825 76.090 88.225 76.490 ;
        RECT 89.825 76.090 90.225 76.490 ;
        RECT 91.825 76.090 92.225 76.490 ;
        RECT 93.825 76.090 94.225 76.490 ;
        RECT 95.825 76.090 96.225 76.490 ;
        RECT 97.825 76.090 98.225 76.490 ;
        RECT 99.825 76.090 100.225 76.490 ;
        RECT 101.825 76.090 102.225 76.490 ;
        RECT 103.825 76.090 104.225 76.490 ;
        RECT 105.825 76.090 106.225 76.490 ;
        RECT 107.825 76.090 108.225 76.490 ;
        RECT 109.825 76.090 110.225 76.490 ;
        RECT 111.825 76.090 112.225 76.490 ;
        RECT 113.825 76.090 114.225 76.490 ;
        RECT 115.825 76.090 116.225 76.490 ;
        RECT 117.825 76.090 118.225 76.490 ;
        RECT 119.825 76.090 120.225 76.490 ;
        RECT 121.825 76.090 122.225 76.490 ;
        RECT 123.825 76.090 124.225 76.490 ;
        RECT 125.825 76.090 126.225 76.490 ;
        RECT 127.825 76.090 128.225 76.490 ;
        RECT 129.825 76.090 130.225 76.490 ;
        RECT 131.825 76.090 132.225 76.490 ;
        RECT 133.825 76.090 134.225 76.490 ;
        RECT 135.825 76.090 136.225 76.490 ;
        RECT 137.825 76.090 138.225 76.490 ;
        RECT 139.825 76.090 140.225 76.490 ;
        RECT 141.825 76.090 142.225 76.490 ;
        RECT 143.825 76.090 144.225 76.490 ;
        RECT 145.825 76.090 146.225 76.490 ;
        RECT 147.825 76.090 148.225 76.490 ;
        RECT 149.825 76.090 150.225 76.490 ;
        RECT 151.825 76.090 152.225 76.490 ;
        RECT 153.825 76.090 154.225 76.490 ;
        RECT 6.890 75.890 8.540 76.090 ;
        RECT 8.890 75.890 22.540 76.090 ;
        RECT 22.890 75.890 38.540 76.090 ;
        RECT 38.890 75.890 46.540 76.090 ;
        RECT 46.890 75.890 50.540 76.090 ;
        RECT 50.890 75.890 52.540 76.090 ;
        RECT 52.890 75.890 54.540 76.090 ;
        RECT 54.890 75.890 74.540 76.090 ;
        RECT 86.575 75.890 106.225 76.090 ;
        RECT 106.575 75.890 108.225 76.090 ;
        RECT 108.575 75.890 110.225 76.090 ;
        RECT 110.575 75.890 114.225 76.090 ;
        RECT 114.575 75.890 122.225 76.090 ;
        RECT 122.575 75.890 138.225 76.090 ;
        RECT 138.575 75.890 152.225 76.090 ;
        RECT 152.575 75.890 154.225 76.090 ;
        RECT 6.890 75.490 7.290 75.890 ;
        RECT 8.890 75.490 9.290 75.890 ;
        RECT 10.890 75.490 11.290 75.890 ;
        RECT 12.890 75.490 13.290 75.890 ;
        RECT 14.890 75.490 15.290 75.890 ;
        RECT 16.890 75.490 17.290 75.890 ;
        RECT 18.890 75.490 19.290 75.890 ;
        RECT 20.890 75.490 21.290 75.890 ;
        RECT 22.890 75.490 23.290 75.890 ;
        RECT 24.890 75.490 25.290 75.890 ;
        RECT 26.890 75.490 27.290 75.890 ;
        RECT 28.890 75.490 29.290 75.890 ;
        RECT 30.890 75.490 31.290 75.890 ;
        RECT 32.890 75.490 33.290 75.890 ;
        RECT 34.890 75.490 35.290 75.890 ;
        RECT 36.890 75.490 37.290 75.890 ;
        RECT 38.890 75.490 39.290 75.890 ;
        RECT 40.890 75.490 41.290 75.890 ;
        RECT 42.890 75.490 43.290 75.890 ;
        RECT 44.890 75.490 45.290 75.890 ;
        RECT 46.890 75.490 47.290 75.890 ;
        RECT 48.890 75.490 49.290 75.890 ;
        RECT 50.890 75.490 51.290 75.890 ;
        RECT 52.890 75.490 53.290 75.890 ;
        RECT 54.890 75.490 55.290 75.890 ;
        RECT 56.890 75.490 57.290 75.890 ;
        RECT 58.890 75.490 59.290 75.890 ;
        RECT 60.890 75.490 61.290 75.890 ;
        RECT 62.890 75.490 63.290 75.890 ;
        RECT 64.890 75.490 65.290 75.890 ;
        RECT 66.890 75.490 67.290 75.890 ;
        RECT 68.890 75.490 69.290 75.890 ;
        RECT 70.890 75.490 71.290 75.890 ;
        RECT 72.890 75.490 73.290 75.890 ;
        RECT 87.825 75.490 88.225 75.890 ;
        RECT 89.825 75.490 90.225 75.890 ;
        RECT 91.825 75.490 92.225 75.890 ;
        RECT 93.825 75.490 94.225 75.890 ;
        RECT 95.825 75.490 96.225 75.890 ;
        RECT 97.825 75.490 98.225 75.890 ;
        RECT 99.825 75.490 100.225 75.890 ;
        RECT 101.825 75.490 102.225 75.890 ;
        RECT 103.825 75.490 104.225 75.890 ;
        RECT 105.825 75.490 106.225 75.890 ;
        RECT 107.825 75.490 108.225 75.890 ;
        RECT 109.825 75.490 110.225 75.890 ;
        RECT 111.825 75.490 112.225 75.890 ;
        RECT 113.825 75.490 114.225 75.890 ;
        RECT 115.825 75.490 116.225 75.890 ;
        RECT 117.825 75.490 118.225 75.890 ;
        RECT 119.825 75.490 120.225 75.890 ;
        RECT 121.825 75.490 122.225 75.890 ;
        RECT 123.825 75.490 124.225 75.890 ;
        RECT 125.825 75.490 126.225 75.890 ;
        RECT 127.825 75.490 128.225 75.890 ;
        RECT 129.825 75.490 130.225 75.890 ;
        RECT 131.825 75.490 132.225 75.890 ;
        RECT 133.825 75.490 134.225 75.890 ;
        RECT 135.825 75.490 136.225 75.890 ;
        RECT 137.825 75.490 138.225 75.890 ;
        RECT 139.825 75.490 140.225 75.890 ;
        RECT 141.825 75.490 142.225 75.890 ;
        RECT 143.825 75.490 144.225 75.890 ;
        RECT 145.825 75.490 146.225 75.890 ;
        RECT 147.825 75.490 148.225 75.890 ;
        RECT 149.825 75.490 150.225 75.890 ;
        RECT 151.825 75.490 152.225 75.890 ;
        RECT 153.825 75.490 154.225 75.890 ;
        RECT 6.960 74.640 7.220 75.490 ;
        RECT 8.990 74.640 9.190 75.490 ;
        RECT 10.990 74.640 11.190 75.490 ;
        RECT 12.990 74.640 13.190 75.490 ;
        RECT 14.990 74.640 15.190 75.490 ;
        RECT 16.990 74.640 17.190 75.490 ;
        RECT 18.990 74.640 19.190 75.490 ;
        RECT 20.990 74.640 21.190 75.490 ;
        RECT 22.990 74.640 23.190 75.490 ;
        RECT 24.990 74.640 25.190 75.490 ;
        RECT 26.990 74.640 27.190 75.490 ;
        RECT 28.990 74.640 29.190 75.490 ;
        RECT 30.990 74.640 31.190 75.490 ;
        RECT 32.990 74.640 33.190 75.490 ;
        RECT 34.990 74.640 35.190 75.490 ;
        RECT 36.990 74.640 37.190 75.490 ;
        RECT 38.990 74.640 39.190 75.490 ;
        RECT 40.990 74.640 41.190 75.490 ;
        RECT 42.990 74.640 43.190 75.490 ;
        RECT 44.990 74.640 45.190 75.490 ;
        RECT 46.990 74.640 47.190 75.490 ;
        RECT 48.990 74.640 49.190 75.490 ;
        RECT 50.990 74.640 51.190 75.490 ;
        RECT 52.990 74.640 53.190 75.490 ;
        RECT 54.990 74.640 55.190 75.490 ;
        RECT 56.990 74.640 57.190 75.490 ;
        RECT 58.990 74.640 59.190 75.490 ;
        RECT 101.925 74.640 102.125 75.490 ;
        RECT 103.925 74.640 104.125 75.490 ;
        RECT 105.925 74.640 106.125 75.490 ;
        RECT 107.925 74.640 108.125 75.490 ;
        RECT 109.925 74.640 110.125 75.490 ;
        RECT 111.925 74.640 112.125 75.490 ;
        RECT 113.925 74.640 114.125 75.490 ;
        RECT 115.925 74.640 116.125 75.490 ;
        RECT 117.925 74.640 118.125 75.490 ;
        RECT 119.925 74.640 120.125 75.490 ;
        RECT 121.925 74.640 122.125 75.490 ;
        RECT 123.925 74.640 124.125 75.490 ;
        RECT 125.925 74.640 126.125 75.490 ;
        RECT 127.925 74.640 128.125 75.490 ;
        RECT 129.925 74.640 130.125 75.490 ;
        RECT 131.925 74.640 132.125 75.490 ;
        RECT 133.925 74.640 134.125 75.490 ;
        RECT 135.925 74.640 136.125 75.490 ;
        RECT 137.925 74.640 138.125 75.490 ;
        RECT 139.925 74.640 140.125 75.490 ;
        RECT 141.925 74.640 142.125 75.490 ;
        RECT 143.925 74.640 144.125 75.490 ;
        RECT 145.925 74.640 146.125 75.490 ;
        RECT 147.925 74.640 148.125 75.490 ;
        RECT 149.925 74.640 150.125 75.490 ;
        RECT 151.925 74.640 152.125 75.490 ;
        RECT 153.895 74.640 154.155 75.490 ;
        RECT 6.890 74.240 7.290 74.640 ;
        RECT 8.890 74.240 9.290 74.640 ;
        RECT 10.890 74.240 11.290 74.640 ;
        RECT 12.890 74.240 13.290 74.640 ;
        RECT 14.890 74.240 15.290 74.640 ;
        RECT 16.890 74.240 17.290 74.640 ;
        RECT 18.890 74.240 19.290 74.640 ;
        RECT 20.890 74.240 21.290 74.640 ;
        RECT 22.890 74.240 23.290 74.640 ;
        RECT 24.890 74.240 25.290 74.640 ;
        RECT 26.890 74.240 27.290 74.640 ;
        RECT 28.890 74.240 29.290 74.640 ;
        RECT 30.890 74.240 31.290 74.640 ;
        RECT 32.890 74.240 33.290 74.640 ;
        RECT 34.890 74.240 35.290 74.640 ;
        RECT 36.890 74.240 37.290 74.640 ;
        RECT 38.890 74.240 39.290 74.640 ;
        RECT 40.890 74.240 41.290 74.640 ;
        RECT 42.890 74.240 43.290 74.640 ;
        RECT 44.890 74.240 45.290 74.640 ;
        RECT 46.890 74.240 47.290 74.640 ;
        RECT 48.890 74.240 49.290 74.640 ;
        RECT 50.890 74.240 51.290 74.640 ;
        RECT 52.890 74.240 53.290 74.640 ;
        RECT 54.890 74.240 55.290 74.640 ;
        RECT 56.890 74.240 57.290 74.640 ;
        RECT 58.890 74.240 59.290 74.640 ;
        RECT 60.890 74.240 61.290 74.640 ;
        RECT 62.890 74.240 63.290 74.640 ;
        RECT 64.890 74.240 65.290 74.640 ;
        RECT 66.890 74.240 67.290 74.640 ;
        RECT 68.890 74.240 69.290 74.640 ;
        RECT 70.890 74.240 71.290 74.640 ;
        RECT 72.890 74.240 73.290 74.640 ;
        RECT 87.825 74.240 88.225 74.640 ;
        RECT 89.825 74.240 90.225 74.640 ;
        RECT 91.825 74.240 92.225 74.640 ;
        RECT 93.825 74.240 94.225 74.640 ;
        RECT 95.825 74.240 96.225 74.640 ;
        RECT 97.825 74.240 98.225 74.640 ;
        RECT 99.825 74.240 100.225 74.640 ;
        RECT 101.825 74.240 102.225 74.640 ;
        RECT 103.825 74.240 104.225 74.640 ;
        RECT 105.825 74.240 106.225 74.640 ;
        RECT 107.825 74.240 108.225 74.640 ;
        RECT 109.825 74.240 110.225 74.640 ;
        RECT 111.825 74.240 112.225 74.640 ;
        RECT 113.825 74.240 114.225 74.640 ;
        RECT 115.825 74.240 116.225 74.640 ;
        RECT 117.825 74.240 118.225 74.640 ;
        RECT 119.825 74.240 120.225 74.640 ;
        RECT 121.825 74.240 122.225 74.640 ;
        RECT 123.825 74.240 124.225 74.640 ;
        RECT 125.825 74.240 126.225 74.640 ;
        RECT 127.825 74.240 128.225 74.640 ;
        RECT 129.825 74.240 130.225 74.640 ;
        RECT 131.825 74.240 132.225 74.640 ;
        RECT 133.825 74.240 134.225 74.640 ;
        RECT 135.825 74.240 136.225 74.640 ;
        RECT 137.825 74.240 138.225 74.640 ;
        RECT 139.825 74.240 140.225 74.640 ;
        RECT 141.825 74.240 142.225 74.640 ;
        RECT 143.825 74.240 144.225 74.640 ;
        RECT 145.825 74.240 146.225 74.640 ;
        RECT 147.825 74.240 148.225 74.640 ;
        RECT 149.825 74.240 150.225 74.640 ;
        RECT 151.825 74.240 152.225 74.640 ;
        RECT 153.825 74.240 154.225 74.640 ;
        RECT 6.890 74.040 8.540 74.240 ;
        RECT 8.890 74.040 22.540 74.240 ;
        RECT 22.890 74.040 38.540 74.240 ;
        RECT 38.890 74.040 46.540 74.240 ;
        RECT 46.890 74.040 50.540 74.240 ;
        RECT 50.890 74.040 52.540 74.240 ;
        RECT 52.890 74.040 54.540 74.240 ;
        RECT 54.890 74.040 60.540 74.240 ;
        RECT 60.890 74.040 74.540 74.240 ;
        RECT 86.575 74.040 100.225 74.240 ;
        RECT 100.575 74.040 106.225 74.240 ;
        RECT 106.575 74.040 108.225 74.240 ;
        RECT 108.575 74.040 110.225 74.240 ;
        RECT 110.575 74.040 114.225 74.240 ;
        RECT 114.575 74.040 122.225 74.240 ;
        RECT 122.575 74.040 138.225 74.240 ;
        RECT 138.575 74.040 152.225 74.240 ;
        RECT 152.575 74.040 154.225 74.240 ;
        RECT 6.890 73.640 7.290 74.040 ;
        RECT 8.890 73.640 9.290 74.040 ;
        RECT 10.890 73.640 11.290 74.040 ;
        RECT 12.890 73.640 13.290 74.040 ;
        RECT 14.890 73.640 15.290 74.040 ;
        RECT 16.890 73.640 17.290 74.040 ;
        RECT 18.890 73.640 19.290 74.040 ;
        RECT 20.890 73.640 21.290 74.040 ;
        RECT 22.890 73.640 23.290 74.040 ;
        RECT 24.890 73.640 25.290 74.040 ;
        RECT 26.890 73.640 27.290 74.040 ;
        RECT 28.890 73.640 29.290 74.040 ;
        RECT 30.890 73.640 31.290 74.040 ;
        RECT 32.890 73.640 33.290 74.040 ;
        RECT 34.890 73.640 35.290 74.040 ;
        RECT 36.890 73.640 37.290 74.040 ;
        RECT 38.890 73.640 39.290 74.040 ;
        RECT 40.890 73.640 41.290 74.040 ;
        RECT 42.890 73.640 43.290 74.040 ;
        RECT 44.890 73.640 45.290 74.040 ;
        RECT 46.890 73.640 47.290 74.040 ;
        RECT 48.890 73.640 49.290 74.040 ;
        RECT 50.890 73.640 51.290 74.040 ;
        RECT 52.890 73.640 53.290 74.040 ;
        RECT 54.890 73.640 55.290 74.040 ;
        RECT 56.890 73.640 57.290 74.040 ;
        RECT 58.890 73.640 59.290 74.040 ;
        RECT 60.890 73.640 61.290 74.040 ;
        RECT 62.890 73.640 63.290 74.040 ;
        RECT 64.890 73.640 65.290 74.040 ;
        RECT 66.890 73.640 67.290 74.040 ;
        RECT 68.890 73.640 69.290 74.040 ;
        RECT 70.890 73.640 71.290 74.040 ;
        RECT 72.890 73.640 73.290 74.040 ;
        RECT 87.825 73.640 88.225 74.040 ;
        RECT 89.825 73.640 90.225 74.040 ;
        RECT 91.825 73.640 92.225 74.040 ;
        RECT 93.825 73.640 94.225 74.040 ;
        RECT 95.825 73.640 96.225 74.040 ;
        RECT 97.825 73.640 98.225 74.040 ;
        RECT 99.825 73.640 100.225 74.040 ;
        RECT 101.825 73.640 102.225 74.040 ;
        RECT 103.825 73.640 104.225 74.040 ;
        RECT 105.825 73.640 106.225 74.040 ;
        RECT 107.825 73.640 108.225 74.040 ;
        RECT 109.825 73.640 110.225 74.040 ;
        RECT 111.825 73.640 112.225 74.040 ;
        RECT 113.825 73.640 114.225 74.040 ;
        RECT 115.825 73.640 116.225 74.040 ;
        RECT 117.825 73.640 118.225 74.040 ;
        RECT 119.825 73.640 120.225 74.040 ;
        RECT 121.825 73.640 122.225 74.040 ;
        RECT 123.825 73.640 124.225 74.040 ;
        RECT 125.825 73.640 126.225 74.040 ;
        RECT 127.825 73.640 128.225 74.040 ;
        RECT 129.825 73.640 130.225 74.040 ;
        RECT 131.825 73.640 132.225 74.040 ;
        RECT 133.825 73.640 134.225 74.040 ;
        RECT 135.825 73.640 136.225 74.040 ;
        RECT 137.825 73.640 138.225 74.040 ;
        RECT 139.825 73.640 140.225 74.040 ;
        RECT 141.825 73.640 142.225 74.040 ;
        RECT 143.825 73.640 144.225 74.040 ;
        RECT 145.825 73.640 146.225 74.040 ;
        RECT 147.825 73.640 148.225 74.040 ;
        RECT 149.825 73.640 150.225 74.040 ;
        RECT 151.825 73.640 152.225 74.040 ;
        RECT 153.825 73.640 154.225 74.040 ;
        RECT 6.960 72.790 7.220 73.640 ;
        RECT 8.990 72.790 9.190 73.640 ;
        RECT 10.990 72.790 11.190 73.640 ;
        RECT 12.990 72.790 13.190 73.640 ;
        RECT 14.990 72.790 15.190 73.640 ;
        RECT 16.990 72.790 17.190 73.640 ;
        RECT 18.990 72.790 19.190 73.640 ;
        RECT 20.990 72.790 21.190 73.640 ;
        RECT 22.990 72.790 23.190 73.640 ;
        RECT 24.990 72.790 25.190 73.640 ;
        RECT 26.990 72.790 27.190 73.640 ;
        RECT 28.990 72.790 29.190 73.640 ;
        RECT 30.990 72.790 31.190 73.640 ;
        RECT 32.990 72.790 33.190 73.640 ;
        RECT 34.990 72.790 35.190 73.640 ;
        RECT 36.990 72.790 37.190 73.640 ;
        RECT 38.990 72.790 39.190 73.640 ;
        RECT 40.990 72.790 41.190 73.640 ;
        RECT 42.990 72.790 43.190 73.640 ;
        RECT 44.990 72.790 45.190 73.640 ;
        RECT 46.990 72.790 47.190 73.640 ;
        RECT 48.990 72.790 49.190 73.640 ;
        RECT 50.990 72.790 51.190 73.640 ;
        RECT 52.990 72.790 53.190 73.640 ;
        RECT 54.990 72.790 55.190 73.640 ;
        RECT 56.990 72.790 57.190 73.640 ;
        RECT 58.990 72.790 59.190 73.640 ;
        RECT 60.990 72.790 61.190 73.640 ;
        RECT 62.990 72.790 63.190 73.640 ;
        RECT 97.925 72.790 98.125 73.640 ;
        RECT 99.925 72.790 100.125 73.640 ;
        RECT 101.925 72.790 102.125 73.640 ;
        RECT 103.925 72.790 104.125 73.640 ;
        RECT 105.925 72.790 106.125 73.640 ;
        RECT 107.925 72.790 108.125 73.640 ;
        RECT 109.925 72.790 110.125 73.640 ;
        RECT 111.925 72.790 112.125 73.640 ;
        RECT 113.925 72.790 114.125 73.640 ;
        RECT 115.925 72.790 116.125 73.640 ;
        RECT 117.925 72.790 118.125 73.640 ;
        RECT 119.925 72.790 120.125 73.640 ;
        RECT 121.925 72.790 122.125 73.640 ;
        RECT 123.925 72.790 124.125 73.640 ;
        RECT 125.925 72.790 126.125 73.640 ;
        RECT 127.925 72.790 128.125 73.640 ;
        RECT 129.925 72.790 130.125 73.640 ;
        RECT 131.925 72.790 132.125 73.640 ;
        RECT 133.925 72.790 134.125 73.640 ;
        RECT 135.925 72.790 136.125 73.640 ;
        RECT 137.925 72.790 138.125 73.640 ;
        RECT 139.925 72.790 140.125 73.640 ;
        RECT 141.925 72.790 142.125 73.640 ;
        RECT 143.925 72.790 144.125 73.640 ;
        RECT 145.925 72.790 146.125 73.640 ;
        RECT 147.925 72.790 148.125 73.640 ;
        RECT 149.925 72.790 150.125 73.640 ;
        RECT 151.925 72.790 152.125 73.640 ;
        RECT 153.895 72.790 154.155 73.640 ;
        RECT 6.890 72.390 7.290 72.790 ;
        RECT 8.890 72.390 9.290 72.790 ;
        RECT 10.890 72.390 11.290 72.790 ;
        RECT 12.890 72.390 13.290 72.790 ;
        RECT 14.890 72.390 15.290 72.790 ;
        RECT 16.890 72.390 17.290 72.790 ;
        RECT 18.890 72.390 19.290 72.790 ;
        RECT 20.890 72.390 21.290 72.790 ;
        RECT 22.890 72.390 23.290 72.790 ;
        RECT 24.890 72.390 25.290 72.790 ;
        RECT 26.890 72.390 27.290 72.790 ;
        RECT 28.890 72.390 29.290 72.790 ;
        RECT 30.890 72.390 31.290 72.790 ;
        RECT 32.890 72.390 33.290 72.790 ;
        RECT 34.890 72.390 35.290 72.790 ;
        RECT 36.890 72.390 37.290 72.790 ;
        RECT 38.890 72.390 39.290 72.790 ;
        RECT 40.890 72.390 41.290 72.790 ;
        RECT 42.890 72.390 43.290 72.790 ;
        RECT 44.890 72.390 45.290 72.790 ;
        RECT 46.890 72.390 47.290 72.790 ;
        RECT 48.890 72.390 49.290 72.790 ;
        RECT 50.890 72.390 51.290 72.790 ;
        RECT 52.890 72.390 53.290 72.790 ;
        RECT 54.890 72.390 55.290 72.790 ;
        RECT 56.890 72.390 57.290 72.790 ;
        RECT 58.890 72.390 59.290 72.790 ;
        RECT 60.890 72.390 61.290 72.790 ;
        RECT 62.890 72.390 63.290 72.790 ;
        RECT 64.890 72.390 65.290 72.790 ;
        RECT 66.890 72.390 67.290 72.790 ;
        RECT 68.890 72.390 69.290 72.790 ;
        RECT 70.890 72.390 71.290 72.790 ;
        RECT 72.890 72.390 73.290 72.790 ;
        RECT 87.825 72.390 88.225 72.790 ;
        RECT 89.825 72.390 90.225 72.790 ;
        RECT 91.825 72.390 92.225 72.790 ;
        RECT 93.825 72.390 94.225 72.790 ;
        RECT 95.825 72.390 96.225 72.790 ;
        RECT 97.825 72.390 98.225 72.790 ;
        RECT 99.825 72.390 100.225 72.790 ;
        RECT 101.825 72.390 102.225 72.790 ;
        RECT 103.825 72.390 104.225 72.790 ;
        RECT 105.825 72.390 106.225 72.790 ;
        RECT 107.825 72.390 108.225 72.790 ;
        RECT 109.825 72.390 110.225 72.790 ;
        RECT 111.825 72.390 112.225 72.790 ;
        RECT 113.825 72.390 114.225 72.790 ;
        RECT 115.825 72.390 116.225 72.790 ;
        RECT 117.825 72.390 118.225 72.790 ;
        RECT 119.825 72.390 120.225 72.790 ;
        RECT 121.825 72.390 122.225 72.790 ;
        RECT 123.825 72.390 124.225 72.790 ;
        RECT 125.825 72.390 126.225 72.790 ;
        RECT 127.825 72.390 128.225 72.790 ;
        RECT 129.825 72.390 130.225 72.790 ;
        RECT 131.825 72.390 132.225 72.790 ;
        RECT 133.825 72.390 134.225 72.790 ;
        RECT 135.825 72.390 136.225 72.790 ;
        RECT 137.825 72.390 138.225 72.790 ;
        RECT 139.825 72.390 140.225 72.790 ;
        RECT 141.825 72.390 142.225 72.790 ;
        RECT 143.825 72.390 144.225 72.790 ;
        RECT 145.825 72.390 146.225 72.790 ;
        RECT 147.825 72.390 148.225 72.790 ;
        RECT 149.825 72.390 150.225 72.790 ;
        RECT 151.825 72.390 152.225 72.790 ;
        RECT 153.825 72.390 154.225 72.790 ;
        RECT 6.890 72.190 8.540 72.390 ;
        RECT 8.890 72.190 22.540 72.390 ;
        RECT 22.890 72.190 38.540 72.390 ;
        RECT 38.890 72.190 46.540 72.390 ;
        RECT 46.890 72.190 50.540 72.390 ;
        RECT 50.890 72.190 52.540 72.390 ;
        RECT 52.890 72.190 54.540 72.390 ;
        RECT 54.890 72.190 60.540 72.390 ;
        RECT 60.890 72.190 64.540 72.390 ;
        RECT 64.890 72.190 74.540 72.390 ;
        RECT 86.575 72.190 96.225 72.390 ;
        RECT 96.575 72.190 100.225 72.390 ;
        RECT 100.575 72.190 106.225 72.390 ;
        RECT 106.575 72.190 108.225 72.390 ;
        RECT 108.575 72.190 110.225 72.390 ;
        RECT 110.575 72.190 114.225 72.390 ;
        RECT 114.575 72.190 122.225 72.390 ;
        RECT 122.575 72.190 138.225 72.390 ;
        RECT 138.575 72.190 152.225 72.390 ;
        RECT 152.575 72.190 154.225 72.390 ;
        RECT 6.890 71.790 7.290 72.190 ;
        RECT 8.890 71.790 9.290 72.190 ;
        RECT 10.890 71.790 11.290 72.190 ;
        RECT 12.890 71.790 13.290 72.190 ;
        RECT 14.890 71.790 15.290 72.190 ;
        RECT 16.890 71.790 17.290 72.190 ;
        RECT 18.890 71.790 19.290 72.190 ;
        RECT 20.890 71.790 21.290 72.190 ;
        RECT 22.890 71.790 23.290 72.190 ;
        RECT 24.890 71.790 25.290 72.190 ;
        RECT 26.890 71.790 27.290 72.190 ;
        RECT 28.890 71.790 29.290 72.190 ;
        RECT 30.890 71.790 31.290 72.190 ;
        RECT 32.890 71.790 33.290 72.190 ;
        RECT 34.890 71.790 35.290 72.190 ;
        RECT 36.890 71.790 37.290 72.190 ;
        RECT 38.890 71.790 39.290 72.190 ;
        RECT 40.890 71.790 41.290 72.190 ;
        RECT 42.890 71.790 43.290 72.190 ;
        RECT 44.890 71.790 45.290 72.190 ;
        RECT 46.890 71.790 47.290 72.190 ;
        RECT 48.890 71.790 49.290 72.190 ;
        RECT 50.890 71.790 51.290 72.190 ;
        RECT 52.890 71.790 53.290 72.190 ;
        RECT 54.890 71.790 55.290 72.190 ;
        RECT 56.890 71.790 57.290 72.190 ;
        RECT 58.890 71.790 59.290 72.190 ;
        RECT 60.890 71.790 61.290 72.190 ;
        RECT 62.890 71.790 63.290 72.190 ;
        RECT 64.890 71.790 65.290 72.190 ;
        RECT 66.890 71.790 67.290 72.190 ;
        RECT 68.890 71.790 69.290 72.190 ;
        RECT 70.890 71.790 71.290 72.190 ;
        RECT 72.890 71.790 73.290 72.190 ;
        RECT 87.825 71.790 88.225 72.190 ;
        RECT 89.825 71.790 90.225 72.190 ;
        RECT 91.825 71.790 92.225 72.190 ;
        RECT 93.825 71.790 94.225 72.190 ;
        RECT 95.825 71.790 96.225 72.190 ;
        RECT 97.825 71.790 98.225 72.190 ;
        RECT 99.825 71.790 100.225 72.190 ;
        RECT 101.825 71.790 102.225 72.190 ;
        RECT 103.825 71.790 104.225 72.190 ;
        RECT 105.825 71.790 106.225 72.190 ;
        RECT 107.825 71.790 108.225 72.190 ;
        RECT 109.825 71.790 110.225 72.190 ;
        RECT 111.825 71.790 112.225 72.190 ;
        RECT 113.825 71.790 114.225 72.190 ;
        RECT 115.825 71.790 116.225 72.190 ;
        RECT 117.825 71.790 118.225 72.190 ;
        RECT 119.825 71.790 120.225 72.190 ;
        RECT 121.825 71.790 122.225 72.190 ;
        RECT 123.825 71.790 124.225 72.190 ;
        RECT 125.825 71.790 126.225 72.190 ;
        RECT 127.825 71.790 128.225 72.190 ;
        RECT 129.825 71.790 130.225 72.190 ;
        RECT 131.825 71.790 132.225 72.190 ;
        RECT 133.825 71.790 134.225 72.190 ;
        RECT 135.825 71.790 136.225 72.190 ;
        RECT 137.825 71.790 138.225 72.190 ;
        RECT 139.825 71.790 140.225 72.190 ;
        RECT 141.825 71.790 142.225 72.190 ;
        RECT 143.825 71.790 144.225 72.190 ;
        RECT 145.825 71.790 146.225 72.190 ;
        RECT 147.825 71.790 148.225 72.190 ;
        RECT 149.825 71.790 150.225 72.190 ;
        RECT 151.825 71.790 152.225 72.190 ;
        RECT 153.825 71.790 154.225 72.190 ;
        RECT 6.960 70.940 7.220 71.790 ;
        RECT 8.990 70.940 9.190 71.790 ;
        RECT 10.990 70.940 11.190 71.790 ;
        RECT 12.990 70.940 13.190 71.790 ;
        RECT 14.990 70.940 15.190 71.790 ;
        RECT 16.990 70.940 17.190 71.790 ;
        RECT 18.990 70.940 19.190 71.790 ;
        RECT 20.990 70.940 21.190 71.790 ;
        RECT 22.990 70.940 23.190 71.790 ;
        RECT 24.990 70.940 25.190 71.790 ;
        RECT 26.990 70.940 27.190 71.790 ;
        RECT 28.990 70.940 29.190 71.790 ;
        RECT 30.990 70.940 31.190 71.790 ;
        RECT 32.990 70.940 33.190 71.790 ;
        RECT 34.990 70.940 35.190 71.790 ;
        RECT 36.990 70.940 37.190 71.790 ;
        RECT 38.990 70.940 39.190 71.790 ;
        RECT 40.990 70.940 41.190 71.790 ;
        RECT 42.990 70.940 43.190 71.790 ;
        RECT 44.990 70.940 45.190 71.790 ;
        RECT 46.990 70.940 47.190 71.790 ;
        RECT 48.990 70.940 49.190 71.790 ;
        RECT 50.990 70.940 51.190 71.790 ;
        RECT 52.990 70.940 53.190 71.790 ;
        RECT 54.990 70.940 55.190 71.790 ;
        RECT 56.990 70.940 57.190 71.790 ;
        RECT 58.990 70.940 59.190 71.790 ;
        RECT 60.990 70.940 61.190 71.790 ;
        RECT 62.990 70.940 63.190 71.790 ;
        RECT 64.990 70.940 65.190 71.790 ;
        RECT 95.925 70.940 96.125 71.790 ;
        RECT 97.925 70.940 98.125 71.790 ;
        RECT 99.925 70.940 100.125 71.790 ;
        RECT 101.925 70.940 102.125 71.790 ;
        RECT 103.925 70.940 104.125 71.790 ;
        RECT 105.925 70.940 106.125 71.790 ;
        RECT 107.925 70.940 108.125 71.790 ;
        RECT 109.925 70.940 110.125 71.790 ;
        RECT 111.925 70.940 112.125 71.790 ;
        RECT 113.925 70.940 114.125 71.790 ;
        RECT 115.925 70.940 116.125 71.790 ;
        RECT 117.925 70.940 118.125 71.790 ;
        RECT 119.925 70.940 120.125 71.790 ;
        RECT 121.925 70.940 122.125 71.790 ;
        RECT 123.925 70.940 124.125 71.790 ;
        RECT 125.925 70.940 126.125 71.790 ;
        RECT 127.925 70.940 128.125 71.790 ;
        RECT 129.925 70.940 130.125 71.790 ;
        RECT 131.925 70.940 132.125 71.790 ;
        RECT 133.925 70.940 134.125 71.790 ;
        RECT 135.925 70.940 136.125 71.790 ;
        RECT 137.925 70.940 138.125 71.790 ;
        RECT 139.925 70.940 140.125 71.790 ;
        RECT 141.925 70.940 142.125 71.790 ;
        RECT 143.925 70.940 144.125 71.790 ;
        RECT 145.925 70.940 146.125 71.790 ;
        RECT 147.925 70.940 148.125 71.790 ;
        RECT 149.925 70.940 150.125 71.790 ;
        RECT 151.925 70.940 152.125 71.790 ;
        RECT 153.895 70.940 154.155 71.790 ;
        RECT 6.890 70.540 7.290 70.940 ;
        RECT 8.890 70.540 9.290 70.940 ;
        RECT 10.890 70.540 11.290 70.940 ;
        RECT 12.890 70.540 13.290 70.940 ;
        RECT 14.890 70.540 15.290 70.940 ;
        RECT 16.890 70.540 17.290 70.940 ;
        RECT 18.890 70.540 19.290 70.940 ;
        RECT 20.890 70.540 21.290 70.940 ;
        RECT 22.890 70.540 23.290 70.940 ;
        RECT 24.890 70.540 25.290 70.940 ;
        RECT 26.890 70.540 27.290 70.940 ;
        RECT 28.890 70.540 29.290 70.940 ;
        RECT 30.890 70.540 31.290 70.940 ;
        RECT 32.890 70.540 33.290 70.940 ;
        RECT 34.890 70.540 35.290 70.940 ;
        RECT 36.890 70.540 37.290 70.940 ;
        RECT 38.890 70.540 39.290 70.940 ;
        RECT 40.890 70.540 41.290 70.940 ;
        RECT 42.890 70.540 43.290 70.940 ;
        RECT 44.890 70.540 45.290 70.940 ;
        RECT 46.890 70.540 47.290 70.940 ;
        RECT 48.890 70.540 49.290 70.940 ;
        RECT 50.890 70.540 51.290 70.940 ;
        RECT 52.890 70.540 53.290 70.940 ;
        RECT 54.890 70.540 55.290 70.940 ;
        RECT 56.890 70.540 57.290 70.940 ;
        RECT 58.890 70.540 59.290 70.940 ;
        RECT 60.890 70.540 61.290 70.940 ;
        RECT 62.890 70.540 63.290 70.940 ;
        RECT 64.890 70.540 65.290 70.940 ;
        RECT 66.890 70.540 67.290 70.940 ;
        RECT 68.890 70.540 69.290 70.940 ;
        RECT 70.890 70.540 71.290 70.940 ;
        RECT 72.890 70.540 73.290 70.940 ;
        RECT 79.880 70.540 80.300 70.620 ;
        RECT 6.890 70.340 8.540 70.540 ;
        RECT 8.890 70.340 22.540 70.540 ;
        RECT 22.890 70.340 38.540 70.540 ;
        RECT 38.890 70.340 46.540 70.540 ;
        RECT 46.890 70.340 50.540 70.540 ;
        RECT 50.890 70.340 52.540 70.540 ;
        RECT 52.890 70.340 54.540 70.540 ;
        RECT 54.890 70.340 60.540 70.540 ;
        RECT 60.890 70.340 64.540 70.540 ;
        RECT 64.890 70.340 66.540 70.540 ;
        RECT 66.890 70.340 80.300 70.540 ;
        RECT 6.890 69.940 7.290 70.340 ;
        RECT 8.890 69.940 9.290 70.340 ;
        RECT 10.890 69.940 11.290 70.340 ;
        RECT 12.890 69.940 13.290 70.340 ;
        RECT 14.890 69.940 15.290 70.340 ;
        RECT 16.890 69.940 17.290 70.340 ;
        RECT 18.890 69.940 19.290 70.340 ;
        RECT 20.890 69.940 21.290 70.340 ;
        RECT 22.890 69.940 23.290 70.340 ;
        RECT 24.890 69.940 25.290 70.340 ;
        RECT 26.890 69.940 27.290 70.340 ;
        RECT 28.890 69.940 29.290 70.340 ;
        RECT 30.890 69.940 31.290 70.340 ;
        RECT 32.890 69.940 33.290 70.340 ;
        RECT 34.890 69.940 35.290 70.340 ;
        RECT 36.890 69.940 37.290 70.340 ;
        RECT 38.890 69.940 39.290 70.340 ;
        RECT 40.890 69.940 41.290 70.340 ;
        RECT 42.890 69.940 43.290 70.340 ;
        RECT 44.890 69.940 45.290 70.340 ;
        RECT 46.890 69.940 47.290 70.340 ;
        RECT 48.890 69.940 49.290 70.340 ;
        RECT 50.890 69.940 51.290 70.340 ;
        RECT 52.890 69.940 53.290 70.340 ;
        RECT 54.890 69.940 55.290 70.340 ;
        RECT 56.890 69.940 57.290 70.340 ;
        RECT 58.890 69.940 59.290 70.340 ;
        RECT 60.890 69.940 61.290 70.340 ;
        RECT 62.890 69.940 63.290 70.340 ;
        RECT 64.890 69.940 65.290 70.340 ;
        RECT 66.890 69.940 67.290 70.340 ;
        RECT 68.890 69.940 69.290 70.340 ;
        RECT 70.890 69.940 71.290 70.340 ;
        RECT 72.890 69.940 73.290 70.340 ;
        RECT 79.880 70.260 80.300 70.340 ;
        RECT 80.815 70.540 81.235 70.620 ;
        RECT 87.825 70.540 88.225 70.940 ;
        RECT 89.825 70.540 90.225 70.940 ;
        RECT 91.825 70.540 92.225 70.940 ;
        RECT 93.825 70.540 94.225 70.940 ;
        RECT 95.825 70.540 96.225 70.940 ;
        RECT 97.825 70.540 98.225 70.940 ;
        RECT 99.825 70.540 100.225 70.940 ;
        RECT 101.825 70.540 102.225 70.940 ;
        RECT 103.825 70.540 104.225 70.940 ;
        RECT 105.825 70.540 106.225 70.940 ;
        RECT 107.825 70.540 108.225 70.940 ;
        RECT 109.825 70.540 110.225 70.940 ;
        RECT 111.825 70.540 112.225 70.940 ;
        RECT 113.825 70.540 114.225 70.940 ;
        RECT 115.825 70.540 116.225 70.940 ;
        RECT 117.825 70.540 118.225 70.940 ;
        RECT 119.825 70.540 120.225 70.940 ;
        RECT 121.825 70.540 122.225 70.940 ;
        RECT 123.825 70.540 124.225 70.940 ;
        RECT 125.825 70.540 126.225 70.940 ;
        RECT 127.825 70.540 128.225 70.940 ;
        RECT 129.825 70.540 130.225 70.940 ;
        RECT 131.825 70.540 132.225 70.940 ;
        RECT 133.825 70.540 134.225 70.940 ;
        RECT 135.825 70.540 136.225 70.940 ;
        RECT 137.825 70.540 138.225 70.940 ;
        RECT 139.825 70.540 140.225 70.940 ;
        RECT 141.825 70.540 142.225 70.940 ;
        RECT 143.825 70.540 144.225 70.940 ;
        RECT 145.825 70.540 146.225 70.940 ;
        RECT 147.825 70.540 148.225 70.940 ;
        RECT 149.825 70.540 150.225 70.940 ;
        RECT 151.825 70.540 152.225 70.940 ;
        RECT 153.825 70.540 154.225 70.940 ;
        RECT 80.815 70.340 94.225 70.540 ;
        RECT 94.575 70.340 96.225 70.540 ;
        RECT 96.575 70.340 100.225 70.540 ;
        RECT 100.575 70.340 106.225 70.540 ;
        RECT 106.575 70.340 108.225 70.540 ;
        RECT 108.575 70.340 110.225 70.540 ;
        RECT 110.575 70.340 114.225 70.540 ;
        RECT 114.575 70.340 122.225 70.540 ;
        RECT 122.575 70.340 138.225 70.540 ;
        RECT 138.575 70.340 152.225 70.540 ;
        RECT 152.575 70.340 154.225 70.540 ;
        RECT 80.815 70.260 81.235 70.340 ;
        RECT 87.825 69.940 88.225 70.340 ;
        RECT 89.825 69.940 90.225 70.340 ;
        RECT 91.825 69.940 92.225 70.340 ;
        RECT 93.825 69.940 94.225 70.340 ;
        RECT 95.825 69.940 96.225 70.340 ;
        RECT 97.825 69.940 98.225 70.340 ;
        RECT 99.825 69.940 100.225 70.340 ;
        RECT 101.825 69.940 102.225 70.340 ;
        RECT 103.825 69.940 104.225 70.340 ;
        RECT 105.825 69.940 106.225 70.340 ;
        RECT 107.825 69.940 108.225 70.340 ;
        RECT 109.825 69.940 110.225 70.340 ;
        RECT 111.825 69.940 112.225 70.340 ;
        RECT 113.825 69.940 114.225 70.340 ;
        RECT 115.825 69.940 116.225 70.340 ;
        RECT 117.825 69.940 118.225 70.340 ;
        RECT 119.825 69.940 120.225 70.340 ;
        RECT 121.825 69.940 122.225 70.340 ;
        RECT 123.825 69.940 124.225 70.340 ;
        RECT 125.825 69.940 126.225 70.340 ;
        RECT 127.825 69.940 128.225 70.340 ;
        RECT 129.825 69.940 130.225 70.340 ;
        RECT 131.825 69.940 132.225 70.340 ;
        RECT 133.825 69.940 134.225 70.340 ;
        RECT 135.825 69.940 136.225 70.340 ;
        RECT 137.825 69.940 138.225 70.340 ;
        RECT 139.825 69.940 140.225 70.340 ;
        RECT 141.825 69.940 142.225 70.340 ;
        RECT 143.825 69.940 144.225 70.340 ;
        RECT 145.825 69.940 146.225 70.340 ;
        RECT 147.825 69.940 148.225 70.340 ;
        RECT 149.825 69.940 150.225 70.340 ;
        RECT 151.825 69.940 152.225 70.340 ;
        RECT 153.825 69.940 154.225 70.340 ;
        RECT 6.960 69.090 7.220 69.940 ;
        RECT 8.990 69.090 9.190 69.940 ;
        RECT 10.990 69.090 11.190 69.940 ;
        RECT 12.990 69.090 13.190 69.940 ;
        RECT 14.990 69.090 15.190 69.940 ;
        RECT 16.990 69.090 17.190 69.940 ;
        RECT 18.990 69.090 19.190 69.940 ;
        RECT 20.990 69.090 21.190 69.940 ;
        RECT 22.990 69.090 23.190 69.940 ;
        RECT 24.990 69.090 25.190 69.940 ;
        RECT 26.990 69.090 27.190 69.940 ;
        RECT 28.990 69.090 29.190 69.940 ;
        RECT 30.990 69.090 31.190 69.940 ;
        RECT 32.990 69.090 33.190 69.940 ;
        RECT 34.990 69.090 35.190 69.940 ;
        RECT 36.990 69.090 37.190 69.940 ;
        RECT 38.990 69.090 39.190 69.940 ;
        RECT 40.990 69.090 41.190 69.940 ;
        RECT 42.990 69.090 43.190 69.940 ;
        RECT 44.990 69.090 45.190 69.940 ;
        RECT 46.990 69.090 47.190 69.940 ;
        RECT 48.990 69.090 49.190 69.940 ;
        RECT 50.990 69.090 51.190 69.940 ;
        RECT 52.990 69.090 53.190 69.940 ;
        RECT 54.990 69.090 55.190 69.940 ;
        RECT 56.990 69.090 57.190 69.940 ;
        RECT 60.990 69.090 61.190 69.940 ;
        RECT 62.990 69.090 63.190 69.940 ;
        RECT 64.990 69.090 65.190 69.940 ;
        RECT 66.990 69.090 67.190 69.940 ;
        RECT 93.925 69.090 94.125 69.940 ;
        RECT 95.925 69.090 96.125 69.940 ;
        RECT 97.925 69.090 98.125 69.940 ;
        RECT 99.925 69.090 100.125 69.940 ;
        RECT 103.925 69.090 104.125 69.940 ;
        RECT 105.925 69.090 106.125 69.940 ;
        RECT 107.925 69.090 108.125 69.940 ;
        RECT 109.925 69.090 110.125 69.940 ;
        RECT 111.925 69.090 112.125 69.940 ;
        RECT 113.925 69.090 114.125 69.940 ;
        RECT 115.925 69.090 116.125 69.940 ;
        RECT 117.925 69.090 118.125 69.940 ;
        RECT 119.925 69.090 120.125 69.940 ;
        RECT 121.925 69.090 122.125 69.940 ;
        RECT 123.925 69.090 124.125 69.940 ;
        RECT 125.925 69.090 126.125 69.940 ;
        RECT 127.925 69.090 128.125 69.940 ;
        RECT 129.925 69.090 130.125 69.940 ;
        RECT 131.925 69.090 132.125 69.940 ;
        RECT 133.925 69.090 134.125 69.940 ;
        RECT 135.925 69.090 136.125 69.940 ;
        RECT 137.925 69.090 138.125 69.940 ;
        RECT 139.925 69.090 140.125 69.940 ;
        RECT 141.925 69.090 142.125 69.940 ;
        RECT 143.925 69.090 144.125 69.940 ;
        RECT 145.925 69.090 146.125 69.940 ;
        RECT 147.925 69.090 148.125 69.940 ;
        RECT 149.925 69.090 150.125 69.940 ;
        RECT 151.925 69.090 152.125 69.940 ;
        RECT 153.895 69.090 154.155 69.940 ;
        RECT 6.890 68.690 7.290 69.090 ;
        RECT 8.890 68.690 9.290 69.090 ;
        RECT 10.890 68.690 11.290 69.090 ;
        RECT 12.890 68.690 13.290 69.090 ;
        RECT 14.890 68.690 15.290 69.090 ;
        RECT 16.890 68.690 17.290 69.090 ;
        RECT 18.890 68.690 19.290 69.090 ;
        RECT 20.890 68.690 21.290 69.090 ;
        RECT 22.890 68.690 23.290 69.090 ;
        RECT 24.890 68.690 25.290 69.090 ;
        RECT 26.890 68.690 27.290 69.090 ;
        RECT 28.890 68.690 29.290 69.090 ;
        RECT 30.890 68.690 31.290 69.090 ;
        RECT 32.890 68.690 33.290 69.090 ;
        RECT 34.890 68.690 35.290 69.090 ;
        RECT 36.890 68.690 37.290 69.090 ;
        RECT 38.890 68.690 39.290 69.090 ;
        RECT 40.890 68.690 41.290 69.090 ;
        RECT 42.890 68.690 43.290 69.090 ;
        RECT 44.890 68.690 45.290 69.090 ;
        RECT 46.890 68.690 47.290 69.090 ;
        RECT 48.890 68.690 49.290 69.090 ;
        RECT 50.890 68.690 51.290 69.090 ;
        RECT 52.890 68.690 53.290 69.090 ;
        RECT 54.890 68.690 55.290 69.090 ;
        RECT 56.890 68.690 57.290 69.090 ;
        RECT 58.890 68.690 59.290 69.090 ;
        RECT 60.890 68.690 61.290 69.090 ;
        RECT 62.890 68.690 63.290 69.090 ;
        RECT 64.890 68.690 65.290 69.090 ;
        RECT 66.890 68.690 67.290 69.090 ;
        RECT 68.890 68.690 69.290 69.090 ;
        RECT 70.890 68.690 71.290 69.090 ;
        RECT 72.890 68.690 73.290 69.090 ;
        RECT 79.430 68.690 79.850 68.770 ;
        RECT 6.890 68.490 8.540 68.690 ;
        RECT 8.890 68.490 22.540 68.690 ;
        RECT 22.890 68.490 38.540 68.690 ;
        RECT 38.890 68.490 46.540 68.690 ;
        RECT 46.890 68.490 50.540 68.690 ;
        RECT 50.890 68.490 52.540 68.690 ;
        RECT 52.890 68.490 54.540 68.690 ;
        RECT 54.890 68.490 58.540 68.690 ;
        RECT 58.890 68.490 64.540 68.690 ;
        RECT 64.890 68.490 66.540 68.690 ;
        RECT 66.890 68.490 68.540 68.690 ;
        RECT 68.890 68.490 79.850 68.690 ;
        RECT 6.890 68.090 7.290 68.490 ;
        RECT 8.890 68.090 9.290 68.490 ;
        RECT 10.890 68.090 11.290 68.490 ;
        RECT 12.890 68.090 13.290 68.490 ;
        RECT 14.890 68.090 15.290 68.490 ;
        RECT 16.890 68.090 17.290 68.490 ;
        RECT 18.890 68.090 19.290 68.490 ;
        RECT 20.890 68.090 21.290 68.490 ;
        RECT 22.890 68.090 23.290 68.490 ;
        RECT 24.890 68.090 25.290 68.490 ;
        RECT 26.890 68.090 27.290 68.490 ;
        RECT 28.890 68.090 29.290 68.490 ;
        RECT 30.890 68.090 31.290 68.490 ;
        RECT 32.890 68.090 33.290 68.490 ;
        RECT 34.890 68.090 35.290 68.490 ;
        RECT 36.890 68.090 37.290 68.490 ;
        RECT 38.890 68.090 39.290 68.490 ;
        RECT 40.890 68.090 41.290 68.490 ;
        RECT 42.890 68.090 43.290 68.490 ;
        RECT 44.890 68.090 45.290 68.490 ;
        RECT 46.890 68.090 47.290 68.490 ;
        RECT 48.890 68.090 49.290 68.490 ;
        RECT 50.890 68.090 51.290 68.490 ;
        RECT 52.890 68.090 53.290 68.490 ;
        RECT 54.890 68.090 55.290 68.490 ;
        RECT 56.890 68.090 57.290 68.490 ;
        RECT 58.890 68.090 59.290 68.490 ;
        RECT 60.890 68.090 61.290 68.490 ;
        RECT 62.890 68.090 63.290 68.490 ;
        RECT 64.890 68.090 65.290 68.490 ;
        RECT 66.890 68.090 67.290 68.490 ;
        RECT 68.890 68.090 69.290 68.490 ;
        RECT 70.890 68.090 71.290 68.490 ;
        RECT 72.890 68.090 73.290 68.490 ;
        RECT 79.430 68.410 79.850 68.490 ;
        RECT 81.265 68.690 81.685 68.770 ;
        RECT 87.825 68.690 88.225 69.090 ;
        RECT 89.825 68.690 90.225 69.090 ;
        RECT 91.825 68.690 92.225 69.090 ;
        RECT 93.825 68.690 94.225 69.090 ;
        RECT 95.825 68.690 96.225 69.090 ;
        RECT 97.825 68.690 98.225 69.090 ;
        RECT 99.825 68.690 100.225 69.090 ;
        RECT 101.825 68.690 102.225 69.090 ;
        RECT 103.825 68.690 104.225 69.090 ;
        RECT 105.825 68.690 106.225 69.090 ;
        RECT 107.825 68.690 108.225 69.090 ;
        RECT 109.825 68.690 110.225 69.090 ;
        RECT 111.825 68.690 112.225 69.090 ;
        RECT 113.825 68.690 114.225 69.090 ;
        RECT 115.825 68.690 116.225 69.090 ;
        RECT 117.825 68.690 118.225 69.090 ;
        RECT 119.825 68.690 120.225 69.090 ;
        RECT 121.825 68.690 122.225 69.090 ;
        RECT 123.825 68.690 124.225 69.090 ;
        RECT 125.825 68.690 126.225 69.090 ;
        RECT 127.825 68.690 128.225 69.090 ;
        RECT 129.825 68.690 130.225 69.090 ;
        RECT 131.825 68.690 132.225 69.090 ;
        RECT 133.825 68.690 134.225 69.090 ;
        RECT 135.825 68.690 136.225 69.090 ;
        RECT 137.825 68.690 138.225 69.090 ;
        RECT 139.825 68.690 140.225 69.090 ;
        RECT 141.825 68.690 142.225 69.090 ;
        RECT 143.825 68.690 144.225 69.090 ;
        RECT 145.825 68.690 146.225 69.090 ;
        RECT 147.825 68.690 148.225 69.090 ;
        RECT 149.825 68.690 150.225 69.090 ;
        RECT 151.825 68.690 152.225 69.090 ;
        RECT 153.825 68.690 154.225 69.090 ;
        RECT 81.265 68.490 92.225 68.690 ;
        RECT 92.575 68.490 94.225 68.690 ;
        RECT 94.575 68.490 96.225 68.690 ;
        RECT 96.575 68.490 102.225 68.690 ;
        RECT 102.575 68.490 106.225 68.690 ;
        RECT 106.575 68.490 108.225 68.690 ;
        RECT 108.575 68.490 110.225 68.690 ;
        RECT 110.575 68.490 114.225 68.690 ;
        RECT 114.575 68.490 122.225 68.690 ;
        RECT 122.575 68.490 138.225 68.690 ;
        RECT 138.575 68.490 152.225 68.690 ;
        RECT 152.575 68.490 154.225 68.690 ;
        RECT 81.265 68.410 81.685 68.490 ;
        RECT 87.825 68.090 88.225 68.490 ;
        RECT 89.825 68.090 90.225 68.490 ;
        RECT 91.825 68.090 92.225 68.490 ;
        RECT 93.825 68.090 94.225 68.490 ;
        RECT 95.825 68.090 96.225 68.490 ;
        RECT 97.825 68.090 98.225 68.490 ;
        RECT 99.825 68.090 100.225 68.490 ;
        RECT 101.825 68.090 102.225 68.490 ;
        RECT 103.825 68.090 104.225 68.490 ;
        RECT 105.825 68.090 106.225 68.490 ;
        RECT 107.825 68.090 108.225 68.490 ;
        RECT 109.825 68.090 110.225 68.490 ;
        RECT 111.825 68.090 112.225 68.490 ;
        RECT 113.825 68.090 114.225 68.490 ;
        RECT 115.825 68.090 116.225 68.490 ;
        RECT 117.825 68.090 118.225 68.490 ;
        RECT 119.825 68.090 120.225 68.490 ;
        RECT 121.825 68.090 122.225 68.490 ;
        RECT 123.825 68.090 124.225 68.490 ;
        RECT 125.825 68.090 126.225 68.490 ;
        RECT 127.825 68.090 128.225 68.490 ;
        RECT 129.825 68.090 130.225 68.490 ;
        RECT 131.825 68.090 132.225 68.490 ;
        RECT 133.825 68.090 134.225 68.490 ;
        RECT 135.825 68.090 136.225 68.490 ;
        RECT 137.825 68.090 138.225 68.490 ;
        RECT 139.825 68.090 140.225 68.490 ;
        RECT 141.825 68.090 142.225 68.490 ;
        RECT 143.825 68.090 144.225 68.490 ;
        RECT 145.825 68.090 146.225 68.490 ;
        RECT 147.825 68.090 148.225 68.490 ;
        RECT 149.825 68.090 150.225 68.490 ;
        RECT 151.825 68.090 152.225 68.490 ;
        RECT 153.825 68.090 154.225 68.490 ;
        RECT 6.960 67.240 7.220 68.090 ;
        RECT 8.990 67.240 9.190 68.090 ;
        RECT 10.990 67.240 11.190 68.090 ;
        RECT 12.990 67.240 13.190 68.090 ;
        RECT 14.990 67.240 15.190 68.090 ;
        RECT 16.990 67.240 17.190 68.090 ;
        RECT 18.990 67.240 19.190 68.090 ;
        RECT 20.990 67.240 21.190 68.090 ;
        RECT 22.990 67.240 23.190 68.090 ;
        RECT 24.990 67.240 25.190 68.090 ;
        RECT 26.990 67.240 27.190 68.090 ;
        RECT 28.990 67.240 29.190 68.090 ;
        RECT 30.990 67.240 31.190 68.090 ;
        RECT 32.990 67.240 33.190 68.090 ;
        RECT 34.990 67.240 35.190 68.090 ;
        RECT 38.990 67.240 39.190 68.090 ;
        RECT 40.990 67.240 41.190 68.090 ;
        RECT 42.990 67.240 43.190 68.090 ;
        RECT 44.990 67.240 45.190 68.090 ;
        RECT 46.990 67.240 47.190 68.090 ;
        RECT 48.990 67.240 49.190 68.090 ;
        RECT 50.990 67.240 51.190 68.090 ;
        RECT 54.990 67.240 55.190 68.090 ;
        RECT 56.990 67.240 57.190 68.090 ;
        RECT 58.990 67.240 59.190 68.090 ;
        RECT 60.990 67.240 61.190 68.090 ;
        RECT 62.990 67.240 63.190 68.090 ;
        RECT 64.990 67.240 65.190 68.090 ;
        RECT 66.990 67.240 67.190 68.090 ;
        RECT 93.925 67.240 94.125 68.090 ;
        RECT 95.925 67.240 96.125 68.090 ;
        RECT 97.925 67.240 98.125 68.090 ;
        RECT 99.925 67.240 100.125 68.090 ;
        RECT 101.925 67.240 102.125 68.090 ;
        RECT 103.925 67.240 104.125 68.090 ;
        RECT 105.925 67.240 106.125 68.090 ;
        RECT 109.925 67.240 110.125 68.090 ;
        RECT 111.925 67.240 112.125 68.090 ;
        RECT 113.925 67.240 114.125 68.090 ;
        RECT 115.925 67.240 116.125 68.090 ;
        RECT 117.925 67.240 118.125 68.090 ;
        RECT 119.925 67.240 120.125 68.090 ;
        RECT 121.925 67.240 122.125 68.090 ;
        RECT 125.925 67.240 126.125 68.090 ;
        RECT 127.925 67.240 128.125 68.090 ;
        RECT 129.925 67.240 130.125 68.090 ;
        RECT 131.925 67.240 132.125 68.090 ;
        RECT 133.925 67.240 134.125 68.090 ;
        RECT 135.925 67.240 136.125 68.090 ;
        RECT 137.925 67.240 138.125 68.090 ;
        RECT 139.925 67.240 140.125 68.090 ;
        RECT 141.925 67.240 142.125 68.090 ;
        RECT 143.925 67.240 144.125 68.090 ;
        RECT 145.925 67.240 146.125 68.090 ;
        RECT 147.925 67.240 148.125 68.090 ;
        RECT 149.925 67.240 150.125 68.090 ;
        RECT 151.925 67.240 152.125 68.090 ;
        RECT 153.895 67.240 154.155 68.090 ;
        RECT 6.890 66.840 7.290 67.240 ;
        RECT 8.890 66.840 9.290 67.240 ;
        RECT 10.890 66.840 11.290 67.240 ;
        RECT 12.890 66.840 13.290 67.240 ;
        RECT 14.890 66.840 15.290 67.240 ;
        RECT 16.890 66.840 17.290 67.240 ;
        RECT 18.890 66.840 19.290 67.240 ;
        RECT 20.890 66.840 21.290 67.240 ;
        RECT 22.890 66.840 23.290 67.240 ;
        RECT 24.890 66.840 25.290 67.240 ;
        RECT 26.890 66.840 27.290 67.240 ;
        RECT 28.890 66.840 29.290 67.240 ;
        RECT 30.890 66.840 31.290 67.240 ;
        RECT 32.890 66.840 33.290 67.240 ;
        RECT 34.890 66.840 35.290 67.240 ;
        RECT 36.890 66.840 37.290 67.240 ;
        RECT 38.890 66.840 39.290 67.240 ;
        RECT 40.890 66.840 41.290 67.240 ;
        RECT 42.890 66.840 43.290 67.240 ;
        RECT 44.890 66.840 45.290 67.240 ;
        RECT 46.890 66.840 47.290 67.240 ;
        RECT 48.890 66.840 49.290 67.240 ;
        RECT 50.890 66.840 51.290 67.240 ;
        RECT 52.890 66.840 53.290 67.240 ;
        RECT 54.890 66.840 55.290 67.240 ;
        RECT 56.890 66.840 57.290 67.240 ;
        RECT 58.890 66.840 59.290 67.240 ;
        RECT 60.890 66.840 61.290 67.240 ;
        RECT 62.890 66.840 63.290 67.240 ;
        RECT 64.890 66.840 65.290 67.240 ;
        RECT 66.890 66.840 67.290 67.240 ;
        RECT 68.890 66.840 69.290 67.240 ;
        RECT 70.890 66.840 71.290 67.240 ;
        RECT 72.890 66.840 73.290 67.240 ;
        RECT 78.980 66.840 79.400 66.920 ;
        RECT 6.890 66.640 8.540 66.840 ;
        RECT 8.890 66.640 22.540 66.840 ;
        RECT 22.890 66.640 36.540 66.840 ;
        RECT 36.890 66.640 46.540 66.840 ;
        RECT 46.890 66.640 50.540 66.840 ;
        RECT 50.890 66.640 52.540 66.840 ;
        RECT 52.890 66.640 58.540 66.840 ;
        RECT 58.890 66.640 64.540 66.840 ;
        RECT 64.890 66.640 66.540 66.840 ;
        RECT 66.890 66.640 68.540 66.840 ;
        RECT 68.890 66.640 70.540 66.840 ;
        RECT 70.890 66.640 79.400 66.840 ;
        RECT 6.890 66.240 7.290 66.640 ;
        RECT 8.890 66.240 9.290 66.640 ;
        RECT 10.890 66.240 11.290 66.640 ;
        RECT 12.890 66.240 13.290 66.640 ;
        RECT 14.890 66.240 15.290 66.640 ;
        RECT 16.890 66.240 17.290 66.640 ;
        RECT 18.890 66.240 19.290 66.640 ;
        RECT 20.890 66.240 21.290 66.640 ;
        RECT 22.890 66.240 23.290 66.640 ;
        RECT 24.890 66.240 25.290 66.640 ;
        RECT 26.890 66.240 27.290 66.640 ;
        RECT 28.890 66.240 29.290 66.640 ;
        RECT 30.890 66.240 31.290 66.640 ;
        RECT 32.890 66.240 33.290 66.640 ;
        RECT 34.890 66.240 35.290 66.640 ;
        RECT 36.890 66.240 37.290 66.640 ;
        RECT 38.890 66.240 39.290 66.640 ;
        RECT 40.890 66.240 41.290 66.640 ;
        RECT 42.890 66.240 43.290 66.640 ;
        RECT 44.890 66.240 45.290 66.640 ;
        RECT 46.890 66.240 47.290 66.640 ;
        RECT 48.890 66.240 49.290 66.640 ;
        RECT 50.890 66.240 51.290 66.640 ;
        RECT 52.890 66.240 53.290 66.640 ;
        RECT 54.890 66.240 55.290 66.640 ;
        RECT 56.890 66.240 57.290 66.640 ;
        RECT 58.890 66.240 59.290 66.640 ;
        RECT 60.890 66.240 61.290 66.640 ;
        RECT 62.890 66.240 63.290 66.640 ;
        RECT 64.890 66.240 65.290 66.640 ;
        RECT 66.890 66.240 67.290 66.640 ;
        RECT 68.890 66.240 69.290 66.640 ;
        RECT 70.890 66.240 71.290 66.640 ;
        RECT 72.890 66.240 73.290 66.640 ;
        RECT 78.980 66.560 79.400 66.640 ;
        RECT 81.715 66.840 82.135 66.920 ;
        RECT 87.825 66.840 88.225 67.240 ;
        RECT 89.825 66.840 90.225 67.240 ;
        RECT 91.825 66.840 92.225 67.240 ;
        RECT 93.825 66.840 94.225 67.240 ;
        RECT 95.825 66.840 96.225 67.240 ;
        RECT 97.825 66.840 98.225 67.240 ;
        RECT 99.825 66.840 100.225 67.240 ;
        RECT 101.825 66.840 102.225 67.240 ;
        RECT 103.825 66.840 104.225 67.240 ;
        RECT 105.825 66.840 106.225 67.240 ;
        RECT 107.825 66.840 108.225 67.240 ;
        RECT 109.825 66.840 110.225 67.240 ;
        RECT 111.825 66.840 112.225 67.240 ;
        RECT 113.825 66.840 114.225 67.240 ;
        RECT 115.825 66.840 116.225 67.240 ;
        RECT 117.825 66.840 118.225 67.240 ;
        RECT 119.825 66.840 120.225 67.240 ;
        RECT 121.825 66.840 122.225 67.240 ;
        RECT 123.825 66.840 124.225 67.240 ;
        RECT 125.825 66.840 126.225 67.240 ;
        RECT 127.825 66.840 128.225 67.240 ;
        RECT 129.825 66.840 130.225 67.240 ;
        RECT 131.825 66.840 132.225 67.240 ;
        RECT 133.825 66.840 134.225 67.240 ;
        RECT 135.825 66.840 136.225 67.240 ;
        RECT 137.825 66.840 138.225 67.240 ;
        RECT 139.825 66.840 140.225 67.240 ;
        RECT 141.825 66.840 142.225 67.240 ;
        RECT 143.825 66.840 144.225 67.240 ;
        RECT 145.825 66.840 146.225 67.240 ;
        RECT 147.825 66.840 148.225 67.240 ;
        RECT 149.825 66.840 150.225 67.240 ;
        RECT 151.825 66.840 152.225 67.240 ;
        RECT 153.825 66.840 154.225 67.240 ;
        RECT 81.715 66.640 90.225 66.840 ;
        RECT 90.575 66.640 92.225 66.840 ;
        RECT 92.575 66.640 94.225 66.840 ;
        RECT 94.575 66.640 96.225 66.840 ;
        RECT 96.575 66.640 102.225 66.840 ;
        RECT 102.575 66.640 108.225 66.840 ;
        RECT 108.575 66.640 110.225 66.840 ;
        RECT 110.575 66.640 114.225 66.840 ;
        RECT 114.575 66.640 124.225 66.840 ;
        RECT 124.575 66.640 138.225 66.840 ;
        RECT 138.575 66.640 152.225 66.840 ;
        RECT 152.575 66.640 154.225 66.840 ;
        RECT 81.715 66.560 82.135 66.640 ;
        RECT 87.825 66.240 88.225 66.640 ;
        RECT 89.825 66.240 90.225 66.640 ;
        RECT 91.825 66.240 92.225 66.640 ;
        RECT 93.825 66.240 94.225 66.640 ;
        RECT 95.825 66.240 96.225 66.640 ;
        RECT 97.825 66.240 98.225 66.640 ;
        RECT 99.825 66.240 100.225 66.640 ;
        RECT 101.825 66.240 102.225 66.640 ;
        RECT 103.825 66.240 104.225 66.640 ;
        RECT 105.825 66.240 106.225 66.640 ;
        RECT 107.825 66.240 108.225 66.640 ;
        RECT 109.825 66.240 110.225 66.640 ;
        RECT 111.825 66.240 112.225 66.640 ;
        RECT 113.825 66.240 114.225 66.640 ;
        RECT 115.825 66.240 116.225 66.640 ;
        RECT 117.825 66.240 118.225 66.640 ;
        RECT 119.825 66.240 120.225 66.640 ;
        RECT 121.825 66.240 122.225 66.640 ;
        RECT 123.825 66.240 124.225 66.640 ;
        RECT 125.825 66.240 126.225 66.640 ;
        RECT 127.825 66.240 128.225 66.640 ;
        RECT 129.825 66.240 130.225 66.640 ;
        RECT 131.825 66.240 132.225 66.640 ;
        RECT 133.825 66.240 134.225 66.640 ;
        RECT 135.825 66.240 136.225 66.640 ;
        RECT 137.825 66.240 138.225 66.640 ;
        RECT 139.825 66.240 140.225 66.640 ;
        RECT 141.825 66.240 142.225 66.640 ;
        RECT 143.825 66.240 144.225 66.640 ;
        RECT 145.825 66.240 146.225 66.640 ;
        RECT 147.825 66.240 148.225 66.640 ;
        RECT 149.825 66.240 150.225 66.640 ;
        RECT 151.825 66.240 152.225 66.640 ;
        RECT 153.825 66.240 154.225 66.640 ;
        RECT 6.960 65.390 7.220 66.240 ;
        RECT 8.990 65.390 9.190 66.240 ;
        RECT 10.990 65.390 11.190 66.240 ;
        RECT 12.990 65.390 13.190 66.240 ;
        RECT 14.990 65.390 15.190 66.240 ;
        RECT 16.990 65.390 17.190 66.240 ;
        RECT 18.990 65.390 19.190 66.240 ;
        RECT 20.990 65.390 21.190 66.240 ;
        RECT 22.990 65.390 23.190 66.240 ;
        RECT 24.990 65.390 25.190 66.240 ;
        RECT 26.990 65.390 27.190 66.240 ;
        RECT 28.990 65.390 29.190 66.240 ;
        RECT 30.990 65.390 31.190 66.240 ;
        RECT 32.990 65.390 33.190 66.240 ;
        RECT 34.990 65.390 35.190 66.240 ;
        RECT 36.990 65.390 37.190 66.240 ;
        RECT 38.990 65.390 39.190 66.240 ;
        RECT 40.990 65.390 41.190 66.240 ;
        RECT 42.990 65.390 43.190 66.240 ;
        RECT 44.990 65.390 45.190 66.240 ;
        RECT 46.990 65.390 47.190 66.240 ;
        RECT 48.990 65.390 49.190 66.240 ;
        RECT 50.990 65.390 51.190 66.240 ;
        RECT 52.990 65.390 53.190 66.240 ;
        RECT 54.990 65.390 55.190 66.240 ;
        RECT 56.990 65.390 57.190 66.240 ;
        RECT 58.990 65.390 59.190 66.240 ;
        RECT 60.990 65.390 61.190 66.240 ;
        RECT 62.990 65.390 63.190 66.240 ;
        RECT 64.990 65.390 65.190 66.240 ;
        RECT 66.990 65.390 67.190 66.240 ;
        RECT 68.990 65.390 69.190 66.240 ;
        RECT 91.925 65.390 92.125 66.240 ;
        RECT 93.925 65.390 94.125 66.240 ;
        RECT 95.925 65.390 96.125 66.240 ;
        RECT 97.925 65.390 98.125 66.240 ;
        RECT 99.925 65.390 100.125 66.240 ;
        RECT 101.925 65.390 102.125 66.240 ;
        RECT 103.925 65.390 104.125 66.240 ;
        RECT 105.925 65.390 106.125 66.240 ;
        RECT 107.925 65.390 108.125 66.240 ;
        RECT 109.925 65.390 110.125 66.240 ;
        RECT 111.925 65.390 112.125 66.240 ;
        RECT 113.925 65.390 114.125 66.240 ;
        RECT 115.925 65.390 116.125 66.240 ;
        RECT 117.925 65.390 118.125 66.240 ;
        RECT 119.925 65.390 120.125 66.240 ;
        RECT 121.925 65.390 122.125 66.240 ;
        RECT 123.925 65.390 124.125 66.240 ;
        RECT 125.925 65.390 126.125 66.240 ;
        RECT 127.925 65.390 128.125 66.240 ;
        RECT 129.925 65.390 130.125 66.240 ;
        RECT 131.925 65.390 132.125 66.240 ;
        RECT 133.925 65.390 134.125 66.240 ;
        RECT 135.925 65.390 136.125 66.240 ;
        RECT 137.925 65.390 138.125 66.240 ;
        RECT 139.925 65.390 140.125 66.240 ;
        RECT 141.925 65.390 142.125 66.240 ;
        RECT 143.925 65.390 144.125 66.240 ;
        RECT 145.925 65.390 146.125 66.240 ;
        RECT 147.925 65.390 148.125 66.240 ;
        RECT 149.925 65.390 150.125 66.240 ;
        RECT 151.925 65.390 152.125 66.240 ;
        RECT 153.895 65.390 154.155 66.240 ;
        RECT 6.890 64.990 7.290 65.390 ;
        RECT 8.890 64.990 9.290 65.390 ;
        RECT 10.890 64.990 11.290 65.390 ;
        RECT 12.890 64.990 13.290 65.390 ;
        RECT 14.890 64.990 15.290 65.390 ;
        RECT 16.890 64.990 17.290 65.390 ;
        RECT 18.890 64.990 19.290 65.390 ;
        RECT 20.890 64.990 21.290 65.390 ;
        RECT 22.890 64.990 23.290 65.390 ;
        RECT 24.890 64.990 25.290 65.390 ;
        RECT 26.890 64.990 27.290 65.390 ;
        RECT 28.890 64.990 29.290 65.390 ;
        RECT 30.890 64.990 31.290 65.390 ;
        RECT 32.890 64.990 33.290 65.390 ;
        RECT 34.890 64.990 35.290 65.390 ;
        RECT 36.890 64.990 37.290 65.390 ;
        RECT 38.890 64.990 39.290 65.390 ;
        RECT 40.890 64.990 41.290 65.390 ;
        RECT 42.890 64.990 43.290 65.390 ;
        RECT 44.890 64.990 45.290 65.390 ;
        RECT 46.890 64.990 47.290 65.390 ;
        RECT 48.890 64.990 49.290 65.390 ;
        RECT 50.890 64.990 51.290 65.390 ;
        RECT 52.890 64.990 53.290 65.390 ;
        RECT 54.890 64.990 55.290 65.390 ;
        RECT 56.890 64.990 57.290 65.390 ;
        RECT 58.890 64.990 59.290 65.390 ;
        RECT 60.890 64.990 61.290 65.390 ;
        RECT 62.890 64.990 63.290 65.390 ;
        RECT 64.890 64.990 65.290 65.390 ;
        RECT 66.890 64.990 67.290 65.390 ;
        RECT 68.890 64.990 69.290 65.390 ;
        RECT 70.890 64.990 71.290 65.390 ;
        RECT 72.890 64.990 73.290 65.390 ;
        RECT 78.530 64.990 78.950 65.070 ;
        RECT 6.890 64.790 8.540 64.990 ;
        RECT 8.890 64.790 22.540 64.990 ;
        RECT 22.890 64.790 36.540 64.990 ;
        RECT 36.890 64.790 46.540 64.990 ;
        RECT 46.890 64.790 50.540 64.990 ;
        RECT 50.890 64.790 52.540 64.990 ;
        RECT 52.890 64.790 58.540 64.990 ;
        RECT 58.890 64.790 64.540 64.990 ;
        RECT 64.890 64.790 66.540 64.990 ;
        RECT 66.890 64.790 68.540 64.990 ;
        RECT 68.890 64.790 70.540 64.990 ;
        RECT 70.890 64.790 78.950 64.990 ;
        RECT 6.890 64.390 7.290 64.790 ;
        RECT 8.890 64.390 9.290 64.790 ;
        RECT 10.890 64.390 11.290 64.790 ;
        RECT 12.890 64.390 13.290 64.790 ;
        RECT 14.890 64.390 15.290 64.790 ;
        RECT 16.890 64.390 17.290 64.790 ;
        RECT 18.890 64.390 19.290 64.790 ;
        RECT 20.890 64.390 21.290 64.790 ;
        RECT 22.890 64.390 23.290 64.790 ;
        RECT 24.890 64.390 25.290 64.790 ;
        RECT 26.890 64.390 27.290 64.790 ;
        RECT 28.890 64.390 29.290 64.790 ;
        RECT 30.890 64.390 31.290 64.790 ;
        RECT 32.890 64.390 33.290 64.790 ;
        RECT 34.890 64.390 35.290 64.790 ;
        RECT 36.890 64.390 37.290 64.790 ;
        RECT 38.890 64.390 39.290 64.790 ;
        RECT 40.890 64.390 41.290 64.790 ;
        RECT 42.890 64.390 43.290 64.790 ;
        RECT 44.890 64.390 45.290 64.790 ;
        RECT 46.890 64.390 47.290 64.790 ;
        RECT 48.890 64.390 49.290 64.790 ;
        RECT 50.890 64.390 51.290 64.790 ;
        RECT 52.890 64.390 53.290 64.790 ;
        RECT 54.890 64.390 55.290 64.790 ;
        RECT 56.890 64.390 57.290 64.790 ;
        RECT 58.890 64.390 59.290 64.790 ;
        RECT 60.890 64.390 61.290 64.790 ;
        RECT 62.890 64.390 63.290 64.790 ;
        RECT 64.890 64.390 65.290 64.790 ;
        RECT 66.890 64.390 67.290 64.790 ;
        RECT 68.890 64.390 69.290 64.790 ;
        RECT 70.890 64.390 71.290 64.790 ;
        RECT 72.890 64.390 73.290 64.790 ;
        RECT 78.530 64.710 78.950 64.790 ;
        RECT 82.165 64.990 82.585 65.070 ;
        RECT 87.825 64.990 88.225 65.390 ;
        RECT 89.825 64.990 90.225 65.390 ;
        RECT 91.825 64.990 92.225 65.390 ;
        RECT 93.825 64.990 94.225 65.390 ;
        RECT 95.825 64.990 96.225 65.390 ;
        RECT 97.825 64.990 98.225 65.390 ;
        RECT 99.825 64.990 100.225 65.390 ;
        RECT 101.825 64.990 102.225 65.390 ;
        RECT 103.825 64.990 104.225 65.390 ;
        RECT 105.825 64.990 106.225 65.390 ;
        RECT 107.825 64.990 108.225 65.390 ;
        RECT 109.825 64.990 110.225 65.390 ;
        RECT 111.825 64.990 112.225 65.390 ;
        RECT 113.825 64.990 114.225 65.390 ;
        RECT 115.825 64.990 116.225 65.390 ;
        RECT 117.825 64.990 118.225 65.390 ;
        RECT 119.825 64.990 120.225 65.390 ;
        RECT 121.825 64.990 122.225 65.390 ;
        RECT 123.825 64.990 124.225 65.390 ;
        RECT 125.825 64.990 126.225 65.390 ;
        RECT 127.825 64.990 128.225 65.390 ;
        RECT 129.825 64.990 130.225 65.390 ;
        RECT 131.825 64.990 132.225 65.390 ;
        RECT 133.825 64.990 134.225 65.390 ;
        RECT 135.825 64.990 136.225 65.390 ;
        RECT 137.825 64.990 138.225 65.390 ;
        RECT 139.825 64.990 140.225 65.390 ;
        RECT 141.825 64.990 142.225 65.390 ;
        RECT 143.825 64.990 144.225 65.390 ;
        RECT 145.825 64.990 146.225 65.390 ;
        RECT 147.825 64.990 148.225 65.390 ;
        RECT 149.825 64.990 150.225 65.390 ;
        RECT 151.825 64.990 152.225 65.390 ;
        RECT 153.825 64.990 154.225 65.390 ;
        RECT 82.165 64.790 90.225 64.990 ;
        RECT 90.575 64.790 92.225 64.990 ;
        RECT 92.575 64.790 94.225 64.990 ;
        RECT 94.575 64.790 96.225 64.990 ;
        RECT 96.575 64.790 102.225 64.990 ;
        RECT 102.575 64.790 108.225 64.990 ;
        RECT 108.575 64.790 110.225 64.990 ;
        RECT 110.575 64.790 114.225 64.990 ;
        RECT 114.575 64.790 124.225 64.990 ;
        RECT 124.575 64.790 138.225 64.990 ;
        RECT 138.575 64.790 152.225 64.990 ;
        RECT 152.575 64.790 154.225 64.990 ;
        RECT 82.165 64.710 82.585 64.790 ;
        RECT 87.825 64.390 88.225 64.790 ;
        RECT 89.825 64.390 90.225 64.790 ;
        RECT 91.825 64.390 92.225 64.790 ;
        RECT 93.825 64.390 94.225 64.790 ;
        RECT 95.825 64.390 96.225 64.790 ;
        RECT 97.825 64.390 98.225 64.790 ;
        RECT 99.825 64.390 100.225 64.790 ;
        RECT 101.825 64.390 102.225 64.790 ;
        RECT 103.825 64.390 104.225 64.790 ;
        RECT 105.825 64.390 106.225 64.790 ;
        RECT 107.825 64.390 108.225 64.790 ;
        RECT 109.825 64.390 110.225 64.790 ;
        RECT 111.825 64.390 112.225 64.790 ;
        RECT 113.825 64.390 114.225 64.790 ;
        RECT 115.825 64.390 116.225 64.790 ;
        RECT 117.825 64.390 118.225 64.790 ;
        RECT 119.825 64.390 120.225 64.790 ;
        RECT 121.825 64.390 122.225 64.790 ;
        RECT 123.825 64.390 124.225 64.790 ;
        RECT 125.825 64.390 126.225 64.790 ;
        RECT 127.825 64.390 128.225 64.790 ;
        RECT 129.825 64.390 130.225 64.790 ;
        RECT 131.825 64.390 132.225 64.790 ;
        RECT 133.825 64.390 134.225 64.790 ;
        RECT 135.825 64.390 136.225 64.790 ;
        RECT 137.825 64.390 138.225 64.790 ;
        RECT 139.825 64.390 140.225 64.790 ;
        RECT 141.825 64.390 142.225 64.790 ;
        RECT 143.825 64.390 144.225 64.790 ;
        RECT 145.825 64.390 146.225 64.790 ;
        RECT 147.825 64.390 148.225 64.790 ;
        RECT 149.825 64.390 150.225 64.790 ;
        RECT 151.825 64.390 152.225 64.790 ;
        RECT 153.825 64.390 154.225 64.790 ;
        RECT 6.960 63.540 7.220 64.390 ;
        RECT 8.990 63.540 9.190 64.390 ;
        RECT 10.990 63.540 11.190 64.390 ;
        RECT 12.990 63.540 13.190 64.390 ;
        RECT 14.990 63.540 15.190 64.390 ;
        RECT 16.990 63.540 17.190 64.390 ;
        RECT 18.990 63.540 19.190 64.390 ;
        RECT 20.990 63.540 21.190 64.390 ;
        RECT 22.990 63.540 23.190 64.390 ;
        RECT 24.990 63.540 25.190 64.390 ;
        RECT 26.990 63.540 27.190 64.390 ;
        RECT 28.990 63.540 29.190 64.390 ;
        RECT 30.990 63.540 31.190 64.390 ;
        RECT 32.990 63.540 33.190 64.390 ;
        RECT 34.990 63.540 35.190 64.390 ;
        RECT 38.990 63.540 39.190 64.390 ;
        RECT 40.990 63.540 41.190 64.390 ;
        RECT 42.990 63.540 43.190 64.390 ;
        RECT 44.990 63.540 45.190 64.390 ;
        RECT 46.990 63.540 47.190 64.390 ;
        RECT 48.990 63.540 49.190 64.390 ;
        RECT 50.990 63.540 51.190 64.390 ;
        RECT 54.990 63.540 55.190 64.390 ;
        RECT 56.990 63.540 57.190 64.390 ;
        RECT 58.990 63.540 59.190 64.390 ;
        RECT 60.990 63.540 61.190 64.390 ;
        RECT 62.990 63.540 63.190 64.390 ;
        RECT 64.990 63.540 65.190 64.390 ;
        RECT 66.990 63.540 67.190 64.390 ;
        RECT 68.990 63.540 69.190 64.390 ;
        RECT 91.925 63.540 92.125 64.390 ;
        RECT 93.925 63.540 94.125 64.390 ;
        RECT 95.925 63.540 96.125 64.390 ;
        RECT 97.925 63.540 98.125 64.390 ;
        RECT 99.925 63.540 100.125 64.390 ;
        RECT 101.925 63.540 102.125 64.390 ;
        RECT 103.925 63.540 104.125 64.390 ;
        RECT 105.925 63.540 106.125 64.390 ;
        RECT 109.925 63.540 110.125 64.390 ;
        RECT 111.925 63.540 112.125 64.390 ;
        RECT 113.925 63.540 114.125 64.390 ;
        RECT 115.925 63.540 116.125 64.390 ;
        RECT 117.925 63.540 118.125 64.390 ;
        RECT 119.925 63.540 120.125 64.390 ;
        RECT 121.925 63.540 122.125 64.390 ;
        RECT 125.925 63.540 126.125 64.390 ;
        RECT 127.925 63.540 128.125 64.390 ;
        RECT 129.925 63.540 130.125 64.390 ;
        RECT 131.925 63.540 132.125 64.390 ;
        RECT 133.925 63.540 134.125 64.390 ;
        RECT 135.925 63.540 136.125 64.390 ;
        RECT 137.925 63.540 138.125 64.390 ;
        RECT 139.925 63.540 140.125 64.390 ;
        RECT 141.925 63.540 142.125 64.390 ;
        RECT 143.925 63.540 144.125 64.390 ;
        RECT 145.925 63.540 146.125 64.390 ;
        RECT 147.925 63.540 148.125 64.390 ;
        RECT 149.925 63.540 150.125 64.390 ;
        RECT 151.925 63.540 152.125 64.390 ;
        RECT 153.895 63.540 154.155 64.390 ;
        RECT 6.890 63.140 7.290 63.540 ;
        RECT 8.890 63.140 9.290 63.540 ;
        RECT 10.890 63.140 11.290 63.540 ;
        RECT 12.890 63.140 13.290 63.540 ;
        RECT 14.890 63.140 15.290 63.540 ;
        RECT 16.890 63.140 17.290 63.540 ;
        RECT 18.890 63.140 19.290 63.540 ;
        RECT 20.890 63.140 21.290 63.540 ;
        RECT 22.890 63.140 23.290 63.540 ;
        RECT 24.890 63.140 25.290 63.540 ;
        RECT 26.890 63.140 27.290 63.540 ;
        RECT 28.890 63.140 29.290 63.540 ;
        RECT 30.890 63.140 31.290 63.540 ;
        RECT 32.890 63.140 33.290 63.540 ;
        RECT 34.890 63.140 35.290 63.540 ;
        RECT 36.890 63.140 37.290 63.540 ;
        RECT 38.890 63.140 39.290 63.540 ;
        RECT 40.890 63.140 41.290 63.540 ;
        RECT 42.890 63.140 43.290 63.540 ;
        RECT 44.890 63.140 45.290 63.540 ;
        RECT 46.890 63.140 47.290 63.540 ;
        RECT 48.890 63.140 49.290 63.540 ;
        RECT 50.890 63.140 51.290 63.540 ;
        RECT 52.890 63.140 53.290 63.540 ;
        RECT 54.890 63.140 55.290 63.540 ;
        RECT 56.890 63.140 57.290 63.540 ;
        RECT 58.890 63.140 59.290 63.540 ;
        RECT 60.890 63.140 61.290 63.540 ;
        RECT 62.890 63.140 63.290 63.540 ;
        RECT 64.890 63.140 65.290 63.540 ;
        RECT 66.890 63.140 67.290 63.540 ;
        RECT 68.890 63.140 69.290 63.540 ;
        RECT 70.890 63.140 71.290 63.540 ;
        RECT 72.890 63.140 73.290 63.540 ;
        RECT 78.080 63.140 78.500 63.220 ;
        RECT 6.890 62.940 8.540 63.140 ;
        RECT 8.890 62.940 22.540 63.140 ;
        RECT 22.890 62.940 38.540 63.140 ;
        RECT 38.890 62.940 46.540 63.140 ;
        RECT 46.890 62.940 50.540 63.140 ;
        RECT 50.890 62.940 52.540 63.140 ;
        RECT 52.890 62.940 54.540 63.140 ;
        RECT 54.890 62.940 58.540 63.140 ;
        RECT 58.890 62.940 64.540 63.140 ;
        RECT 64.890 62.940 66.540 63.140 ;
        RECT 66.890 62.940 68.540 63.140 ;
        RECT 68.890 62.940 78.500 63.140 ;
        RECT 6.890 62.540 7.290 62.940 ;
        RECT 8.890 62.540 9.290 62.940 ;
        RECT 10.890 62.540 11.290 62.940 ;
        RECT 12.890 62.540 13.290 62.940 ;
        RECT 14.890 62.540 15.290 62.940 ;
        RECT 16.890 62.540 17.290 62.940 ;
        RECT 18.890 62.540 19.290 62.940 ;
        RECT 20.890 62.540 21.290 62.940 ;
        RECT 22.890 62.540 23.290 62.940 ;
        RECT 24.890 62.540 25.290 62.940 ;
        RECT 26.890 62.540 27.290 62.940 ;
        RECT 28.890 62.540 29.290 62.940 ;
        RECT 30.890 62.540 31.290 62.940 ;
        RECT 32.890 62.540 33.290 62.940 ;
        RECT 34.890 62.540 35.290 62.940 ;
        RECT 36.890 62.540 37.290 62.940 ;
        RECT 38.890 62.540 39.290 62.940 ;
        RECT 40.890 62.540 41.290 62.940 ;
        RECT 42.890 62.540 43.290 62.940 ;
        RECT 44.890 62.540 45.290 62.940 ;
        RECT 46.890 62.540 47.290 62.940 ;
        RECT 48.890 62.540 49.290 62.940 ;
        RECT 50.890 62.540 51.290 62.940 ;
        RECT 52.890 62.540 53.290 62.940 ;
        RECT 54.890 62.540 55.290 62.940 ;
        RECT 56.890 62.540 57.290 62.940 ;
        RECT 58.890 62.540 59.290 62.940 ;
        RECT 60.890 62.540 61.290 62.940 ;
        RECT 62.890 62.540 63.290 62.940 ;
        RECT 64.890 62.540 65.290 62.940 ;
        RECT 66.890 62.540 67.290 62.940 ;
        RECT 68.890 62.540 69.290 62.940 ;
        RECT 70.890 62.540 71.290 62.940 ;
        RECT 72.890 62.540 73.290 62.940 ;
        RECT 78.080 62.860 78.500 62.940 ;
        RECT 82.615 63.140 83.035 63.220 ;
        RECT 87.825 63.140 88.225 63.540 ;
        RECT 89.825 63.140 90.225 63.540 ;
        RECT 91.825 63.140 92.225 63.540 ;
        RECT 93.825 63.140 94.225 63.540 ;
        RECT 95.825 63.140 96.225 63.540 ;
        RECT 97.825 63.140 98.225 63.540 ;
        RECT 99.825 63.140 100.225 63.540 ;
        RECT 101.825 63.140 102.225 63.540 ;
        RECT 103.825 63.140 104.225 63.540 ;
        RECT 105.825 63.140 106.225 63.540 ;
        RECT 107.825 63.140 108.225 63.540 ;
        RECT 109.825 63.140 110.225 63.540 ;
        RECT 111.825 63.140 112.225 63.540 ;
        RECT 113.825 63.140 114.225 63.540 ;
        RECT 115.825 63.140 116.225 63.540 ;
        RECT 117.825 63.140 118.225 63.540 ;
        RECT 119.825 63.140 120.225 63.540 ;
        RECT 121.825 63.140 122.225 63.540 ;
        RECT 123.825 63.140 124.225 63.540 ;
        RECT 125.825 63.140 126.225 63.540 ;
        RECT 127.825 63.140 128.225 63.540 ;
        RECT 129.825 63.140 130.225 63.540 ;
        RECT 131.825 63.140 132.225 63.540 ;
        RECT 133.825 63.140 134.225 63.540 ;
        RECT 135.825 63.140 136.225 63.540 ;
        RECT 137.825 63.140 138.225 63.540 ;
        RECT 139.825 63.140 140.225 63.540 ;
        RECT 141.825 63.140 142.225 63.540 ;
        RECT 143.825 63.140 144.225 63.540 ;
        RECT 145.825 63.140 146.225 63.540 ;
        RECT 147.825 63.140 148.225 63.540 ;
        RECT 149.825 63.140 150.225 63.540 ;
        RECT 151.825 63.140 152.225 63.540 ;
        RECT 153.825 63.140 154.225 63.540 ;
        RECT 82.615 62.940 92.225 63.140 ;
        RECT 92.575 62.940 94.225 63.140 ;
        RECT 94.575 62.940 96.225 63.140 ;
        RECT 96.575 62.940 102.225 63.140 ;
        RECT 102.575 62.940 106.225 63.140 ;
        RECT 106.575 62.940 108.225 63.140 ;
        RECT 108.575 62.940 110.225 63.140 ;
        RECT 110.575 62.940 114.225 63.140 ;
        RECT 114.575 62.940 122.225 63.140 ;
        RECT 122.575 62.940 138.225 63.140 ;
        RECT 138.575 62.940 152.225 63.140 ;
        RECT 152.575 62.940 154.225 63.140 ;
        RECT 82.615 62.860 83.035 62.940 ;
        RECT 87.825 62.540 88.225 62.940 ;
        RECT 89.825 62.540 90.225 62.940 ;
        RECT 91.825 62.540 92.225 62.940 ;
        RECT 93.825 62.540 94.225 62.940 ;
        RECT 95.825 62.540 96.225 62.940 ;
        RECT 97.825 62.540 98.225 62.940 ;
        RECT 99.825 62.540 100.225 62.940 ;
        RECT 101.825 62.540 102.225 62.940 ;
        RECT 103.825 62.540 104.225 62.940 ;
        RECT 105.825 62.540 106.225 62.940 ;
        RECT 107.825 62.540 108.225 62.940 ;
        RECT 109.825 62.540 110.225 62.940 ;
        RECT 111.825 62.540 112.225 62.940 ;
        RECT 113.825 62.540 114.225 62.940 ;
        RECT 115.825 62.540 116.225 62.940 ;
        RECT 117.825 62.540 118.225 62.940 ;
        RECT 119.825 62.540 120.225 62.940 ;
        RECT 121.825 62.540 122.225 62.940 ;
        RECT 123.825 62.540 124.225 62.940 ;
        RECT 125.825 62.540 126.225 62.940 ;
        RECT 127.825 62.540 128.225 62.940 ;
        RECT 129.825 62.540 130.225 62.940 ;
        RECT 131.825 62.540 132.225 62.940 ;
        RECT 133.825 62.540 134.225 62.940 ;
        RECT 135.825 62.540 136.225 62.940 ;
        RECT 137.825 62.540 138.225 62.940 ;
        RECT 139.825 62.540 140.225 62.940 ;
        RECT 141.825 62.540 142.225 62.940 ;
        RECT 143.825 62.540 144.225 62.940 ;
        RECT 145.825 62.540 146.225 62.940 ;
        RECT 147.825 62.540 148.225 62.940 ;
        RECT 149.825 62.540 150.225 62.940 ;
        RECT 151.825 62.540 152.225 62.940 ;
        RECT 153.825 62.540 154.225 62.940 ;
        RECT 6.960 61.690 7.220 62.540 ;
        RECT 8.990 61.690 9.190 62.540 ;
        RECT 10.990 61.690 11.190 62.540 ;
        RECT 12.990 61.690 13.190 62.540 ;
        RECT 14.990 61.690 15.190 62.540 ;
        RECT 16.990 61.690 17.190 62.540 ;
        RECT 18.990 61.690 19.190 62.540 ;
        RECT 20.990 61.690 21.190 62.540 ;
        RECT 22.990 61.690 23.190 62.540 ;
        RECT 24.990 61.690 25.190 62.540 ;
        RECT 26.990 61.690 27.190 62.540 ;
        RECT 28.990 61.690 29.190 62.540 ;
        RECT 30.990 61.690 31.190 62.540 ;
        RECT 32.990 61.690 33.190 62.540 ;
        RECT 34.990 61.690 35.190 62.540 ;
        RECT 36.990 61.690 37.190 62.540 ;
        RECT 38.990 61.690 39.190 62.540 ;
        RECT 40.990 61.690 41.190 62.540 ;
        RECT 42.990 61.690 43.190 62.540 ;
        RECT 44.990 61.690 45.190 62.540 ;
        RECT 46.990 61.690 47.190 62.540 ;
        RECT 48.990 61.690 49.190 62.540 ;
        RECT 50.990 61.690 51.190 62.540 ;
        RECT 52.990 61.690 53.190 62.540 ;
        RECT 54.990 61.690 55.190 62.540 ;
        RECT 56.990 61.690 57.190 62.540 ;
        RECT 60.990 61.690 61.190 62.540 ;
        RECT 62.990 61.690 63.190 62.540 ;
        RECT 64.990 61.690 65.190 62.540 ;
        RECT 66.990 61.690 67.190 62.540 ;
        RECT 93.925 61.690 94.125 62.540 ;
        RECT 95.925 61.690 96.125 62.540 ;
        RECT 97.925 61.690 98.125 62.540 ;
        RECT 99.925 61.690 100.125 62.540 ;
        RECT 103.925 61.690 104.125 62.540 ;
        RECT 105.925 61.690 106.125 62.540 ;
        RECT 107.925 61.690 108.125 62.540 ;
        RECT 109.925 61.690 110.125 62.540 ;
        RECT 111.925 61.690 112.125 62.540 ;
        RECT 113.925 61.690 114.125 62.540 ;
        RECT 115.925 61.690 116.125 62.540 ;
        RECT 117.925 61.690 118.125 62.540 ;
        RECT 119.925 61.690 120.125 62.540 ;
        RECT 121.925 61.690 122.125 62.540 ;
        RECT 123.925 61.690 124.125 62.540 ;
        RECT 125.925 61.690 126.125 62.540 ;
        RECT 127.925 61.690 128.125 62.540 ;
        RECT 129.925 61.690 130.125 62.540 ;
        RECT 131.925 61.690 132.125 62.540 ;
        RECT 133.925 61.690 134.125 62.540 ;
        RECT 135.925 61.690 136.125 62.540 ;
        RECT 137.925 61.690 138.125 62.540 ;
        RECT 139.925 61.690 140.125 62.540 ;
        RECT 141.925 61.690 142.125 62.540 ;
        RECT 143.925 61.690 144.125 62.540 ;
        RECT 145.925 61.690 146.125 62.540 ;
        RECT 147.925 61.690 148.125 62.540 ;
        RECT 149.925 61.690 150.125 62.540 ;
        RECT 151.925 61.690 152.125 62.540 ;
        RECT 153.895 61.690 154.155 62.540 ;
        RECT 6.890 61.290 7.290 61.690 ;
        RECT 8.890 61.290 9.290 61.690 ;
        RECT 10.890 61.290 11.290 61.690 ;
        RECT 12.890 61.290 13.290 61.690 ;
        RECT 14.890 61.290 15.290 61.690 ;
        RECT 16.890 61.290 17.290 61.690 ;
        RECT 18.890 61.290 19.290 61.690 ;
        RECT 20.890 61.290 21.290 61.690 ;
        RECT 22.890 61.290 23.290 61.690 ;
        RECT 24.890 61.290 25.290 61.690 ;
        RECT 26.890 61.290 27.290 61.690 ;
        RECT 28.890 61.290 29.290 61.690 ;
        RECT 30.890 61.290 31.290 61.690 ;
        RECT 32.890 61.290 33.290 61.690 ;
        RECT 34.890 61.290 35.290 61.690 ;
        RECT 36.890 61.290 37.290 61.690 ;
        RECT 38.890 61.290 39.290 61.690 ;
        RECT 40.890 61.290 41.290 61.690 ;
        RECT 42.890 61.290 43.290 61.690 ;
        RECT 44.890 61.290 45.290 61.690 ;
        RECT 46.890 61.290 47.290 61.690 ;
        RECT 48.890 61.290 49.290 61.690 ;
        RECT 50.890 61.290 51.290 61.690 ;
        RECT 52.890 61.290 53.290 61.690 ;
        RECT 54.890 61.290 55.290 61.690 ;
        RECT 56.890 61.290 57.290 61.690 ;
        RECT 58.890 61.290 59.290 61.690 ;
        RECT 60.890 61.290 61.290 61.690 ;
        RECT 62.890 61.290 63.290 61.690 ;
        RECT 64.890 61.290 65.290 61.690 ;
        RECT 66.890 61.290 67.290 61.690 ;
        RECT 68.890 61.290 69.290 61.690 ;
        RECT 70.890 61.290 71.290 61.690 ;
        RECT 72.890 61.290 73.290 61.690 ;
        RECT 77.630 61.290 78.050 61.370 ;
        RECT 6.890 61.090 8.540 61.290 ;
        RECT 8.890 61.090 22.540 61.290 ;
        RECT 22.890 61.090 38.540 61.290 ;
        RECT 38.890 61.090 46.540 61.290 ;
        RECT 46.890 61.090 50.540 61.290 ;
        RECT 50.890 61.090 52.540 61.290 ;
        RECT 52.890 61.090 54.540 61.290 ;
        RECT 54.890 61.090 60.540 61.290 ;
        RECT 60.890 61.090 64.540 61.290 ;
        RECT 64.890 61.090 66.540 61.290 ;
        RECT 66.890 61.090 68.540 61.290 ;
        RECT 68.890 61.090 78.050 61.290 ;
        RECT 6.890 60.690 7.290 61.090 ;
        RECT 8.890 60.690 9.290 61.090 ;
        RECT 10.890 60.690 11.290 61.090 ;
        RECT 12.890 60.690 13.290 61.090 ;
        RECT 14.890 60.690 15.290 61.090 ;
        RECT 16.890 60.690 17.290 61.090 ;
        RECT 18.890 60.690 19.290 61.090 ;
        RECT 20.890 60.690 21.290 61.090 ;
        RECT 22.890 60.690 23.290 61.090 ;
        RECT 24.890 60.690 25.290 61.090 ;
        RECT 26.890 60.690 27.290 61.090 ;
        RECT 28.890 60.690 29.290 61.090 ;
        RECT 30.890 60.690 31.290 61.090 ;
        RECT 32.890 60.690 33.290 61.090 ;
        RECT 34.890 60.690 35.290 61.090 ;
        RECT 36.890 60.690 37.290 61.090 ;
        RECT 38.890 60.690 39.290 61.090 ;
        RECT 40.890 60.690 41.290 61.090 ;
        RECT 42.890 60.690 43.290 61.090 ;
        RECT 44.890 60.690 45.290 61.090 ;
        RECT 46.890 60.690 47.290 61.090 ;
        RECT 48.890 60.690 49.290 61.090 ;
        RECT 50.890 60.690 51.290 61.090 ;
        RECT 52.890 60.690 53.290 61.090 ;
        RECT 54.890 60.690 55.290 61.090 ;
        RECT 56.890 60.690 57.290 61.090 ;
        RECT 58.890 60.690 59.290 61.090 ;
        RECT 60.890 60.690 61.290 61.090 ;
        RECT 62.890 60.690 63.290 61.090 ;
        RECT 64.890 60.690 65.290 61.090 ;
        RECT 66.890 60.690 67.290 61.090 ;
        RECT 68.890 60.690 69.290 61.090 ;
        RECT 70.890 60.690 71.290 61.090 ;
        RECT 72.890 60.690 73.290 61.090 ;
        RECT 77.630 61.010 78.050 61.090 ;
        RECT 83.065 61.290 83.485 61.370 ;
        RECT 87.825 61.290 88.225 61.690 ;
        RECT 89.825 61.290 90.225 61.690 ;
        RECT 91.825 61.290 92.225 61.690 ;
        RECT 93.825 61.290 94.225 61.690 ;
        RECT 95.825 61.290 96.225 61.690 ;
        RECT 97.825 61.290 98.225 61.690 ;
        RECT 99.825 61.290 100.225 61.690 ;
        RECT 101.825 61.290 102.225 61.690 ;
        RECT 103.825 61.290 104.225 61.690 ;
        RECT 105.825 61.290 106.225 61.690 ;
        RECT 107.825 61.290 108.225 61.690 ;
        RECT 109.825 61.290 110.225 61.690 ;
        RECT 111.825 61.290 112.225 61.690 ;
        RECT 113.825 61.290 114.225 61.690 ;
        RECT 115.825 61.290 116.225 61.690 ;
        RECT 117.825 61.290 118.225 61.690 ;
        RECT 119.825 61.290 120.225 61.690 ;
        RECT 121.825 61.290 122.225 61.690 ;
        RECT 123.825 61.290 124.225 61.690 ;
        RECT 125.825 61.290 126.225 61.690 ;
        RECT 127.825 61.290 128.225 61.690 ;
        RECT 129.825 61.290 130.225 61.690 ;
        RECT 131.825 61.290 132.225 61.690 ;
        RECT 133.825 61.290 134.225 61.690 ;
        RECT 135.825 61.290 136.225 61.690 ;
        RECT 137.825 61.290 138.225 61.690 ;
        RECT 139.825 61.290 140.225 61.690 ;
        RECT 141.825 61.290 142.225 61.690 ;
        RECT 143.825 61.290 144.225 61.690 ;
        RECT 145.825 61.290 146.225 61.690 ;
        RECT 147.825 61.290 148.225 61.690 ;
        RECT 149.825 61.290 150.225 61.690 ;
        RECT 151.825 61.290 152.225 61.690 ;
        RECT 153.825 61.290 154.225 61.690 ;
        RECT 83.065 61.090 92.225 61.290 ;
        RECT 92.575 61.090 94.225 61.290 ;
        RECT 94.575 61.090 96.225 61.290 ;
        RECT 96.575 61.090 100.225 61.290 ;
        RECT 100.575 61.090 106.225 61.290 ;
        RECT 106.575 61.090 108.225 61.290 ;
        RECT 108.575 61.090 110.225 61.290 ;
        RECT 110.575 61.090 114.225 61.290 ;
        RECT 114.575 61.090 122.225 61.290 ;
        RECT 122.575 61.090 138.225 61.290 ;
        RECT 138.575 61.090 152.225 61.290 ;
        RECT 152.575 61.090 154.225 61.290 ;
        RECT 83.065 61.010 83.485 61.090 ;
        RECT 87.825 60.690 88.225 61.090 ;
        RECT 89.825 60.690 90.225 61.090 ;
        RECT 91.825 60.690 92.225 61.090 ;
        RECT 93.825 60.690 94.225 61.090 ;
        RECT 95.825 60.690 96.225 61.090 ;
        RECT 97.825 60.690 98.225 61.090 ;
        RECT 99.825 60.690 100.225 61.090 ;
        RECT 101.825 60.690 102.225 61.090 ;
        RECT 103.825 60.690 104.225 61.090 ;
        RECT 105.825 60.690 106.225 61.090 ;
        RECT 107.825 60.690 108.225 61.090 ;
        RECT 109.825 60.690 110.225 61.090 ;
        RECT 111.825 60.690 112.225 61.090 ;
        RECT 113.825 60.690 114.225 61.090 ;
        RECT 115.825 60.690 116.225 61.090 ;
        RECT 117.825 60.690 118.225 61.090 ;
        RECT 119.825 60.690 120.225 61.090 ;
        RECT 121.825 60.690 122.225 61.090 ;
        RECT 123.825 60.690 124.225 61.090 ;
        RECT 125.825 60.690 126.225 61.090 ;
        RECT 127.825 60.690 128.225 61.090 ;
        RECT 129.825 60.690 130.225 61.090 ;
        RECT 131.825 60.690 132.225 61.090 ;
        RECT 133.825 60.690 134.225 61.090 ;
        RECT 135.825 60.690 136.225 61.090 ;
        RECT 137.825 60.690 138.225 61.090 ;
        RECT 139.825 60.690 140.225 61.090 ;
        RECT 141.825 60.690 142.225 61.090 ;
        RECT 143.825 60.690 144.225 61.090 ;
        RECT 145.825 60.690 146.225 61.090 ;
        RECT 147.825 60.690 148.225 61.090 ;
        RECT 149.825 60.690 150.225 61.090 ;
        RECT 151.825 60.690 152.225 61.090 ;
        RECT 153.825 60.690 154.225 61.090 ;
        RECT 6.960 59.840 7.220 60.690 ;
        RECT 8.990 59.840 9.190 60.690 ;
        RECT 10.990 59.840 11.190 60.690 ;
        RECT 12.990 59.840 13.190 60.690 ;
        RECT 14.990 59.840 15.190 60.690 ;
        RECT 16.990 59.840 17.190 60.690 ;
        RECT 18.990 59.840 19.190 60.690 ;
        RECT 20.990 59.840 21.190 60.690 ;
        RECT 22.990 59.840 23.190 60.690 ;
        RECT 24.990 59.840 25.190 60.690 ;
        RECT 26.990 59.840 27.190 60.690 ;
        RECT 28.990 59.840 29.190 60.690 ;
        RECT 30.990 59.840 31.190 60.690 ;
        RECT 32.990 59.840 33.190 60.690 ;
        RECT 34.990 59.840 35.190 60.690 ;
        RECT 36.990 59.840 37.190 60.690 ;
        RECT 38.990 59.840 39.190 60.690 ;
        RECT 40.990 59.840 41.190 60.690 ;
        RECT 42.990 59.840 43.190 60.690 ;
        RECT 44.990 59.840 45.190 60.690 ;
        RECT 46.990 59.840 47.190 60.690 ;
        RECT 48.990 59.840 49.190 60.690 ;
        RECT 50.990 59.840 51.190 60.690 ;
        RECT 52.990 59.840 53.190 60.690 ;
        RECT 54.990 59.840 55.190 60.690 ;
        RECT 56.990 59.840 57.190 60.690 ;
        RECT 58.990 59.840 59.190 60.690 ;
        RECT 60.990 59.840 61.190 60.690 ;
        RECT 62.990 59.840 63.190 60.690 ;
        RECT 64.990 59.840 65.190 60.690 ;
        RECT 68.990 59.840 69.190 60.690 ;
        RECT 70.990 59.840 71.190 60.690 ;
        RECT 89.925 59.840 90.125 60.690 ;
        RECT 91.925 59.840 92.125 60.690 ;
        RECT 95.925 59.840 96.125 60.690 ;
        RECT 97.925 59.840 98.125 60.690 ;
        RECT 99.925 59.840 100.125 60.690 ;
        RECT 101.925 59.840 102.125 60.690 ;
        RECT 103.925 59.840 104.125 60.690 ;
        RECT 105.925 59.840 106.125 60.690 ;
        RECT 107.925 59.840 108.125 60.690 ;
        RECT 109.925 59.840 110.125 60.690 ;
        RECT 111.925 59.840 112.125 60.690 ;
        RECT 113.925 59.840 114.125 60.690 ;
        RECT 115.925 59.840 116.125 60.690 ;
        RECT 117.925 59.840 118.125 60.690 ;
        RECT 119.925 59.840 120.125 60.690 ;
        RECT 121.925 59.840 122.125 60.690 ;
        RECT 123.925 59.840 124.125 60.690 ;
        RECT 125.925 59.840 126.125 60.690 ;
        RECT 127.925 59.840 128.125 60.690 ;
        RECT 129.925 59.840 130.125 60.690 ;
        RECT 131.925 59.840 132.125 60.690 ;
        RECT 133.925 59.840 134.125 60.690 ;
        RECT 135.925 59.840 136.125 60.690 ;
        RECT 137.925 59.840 138.125 60.690 ;
        RECT 139.925 59.840 140.125 60.690 ;
        RECT 141.925 59.840 142.125 60.690 ;
        RECT 143.925 59.840 144.125 60.690 ;
        RECT 145.925 59.840 146.125 60.690 ;
        RECT 147.925 59.840 148.125 60.690 ;
        RECT 149.925 59.840 150.125 60.690 ;
        RECT 151.925 59.840 152.125 60.690 ;
        RECT 153.895 59.840 154.155 60.690 ;
        RECT 6.890 59.440 7.290 59.840 ;
        RECT 8.890 59.440 9.290 59.840 ;
        RECT 10.890 59.440 11.290 59.840 ;
        RECT 12.890 59.440 13.290 59.840 ;
        RECT 14.890 59.440 15.290 59.840 ;
        RECT 16.890 59.440 17.290 59.840 ;
        RECT 18.890 59.440 19.290 59.840 ;
        RECT 20.890 59.440 21.290 59.840 ;
        RECT 22.890 59.440 23.290 59.840 ;
        RECT 24.890 59.440 25.290 59.840 ;
        RECT 26.890 59.440 27.290 59.840 ;
        RECT 28.890 59.440 29.290 59.840 ;
        RECT 30.890 59.440 31.290 59.840 ;
        RECT 32.890 59.440 33.290 59.840 ;
        RECT 34.890 59.440 35.290 59.840 ;
        RECT 36.890 59.440 37.290 59.840 ;
        RECT 38.890 59.440 39.290 59.840 ;
        RECT 40.890 59.440 41.290 59.840 ;
        RECT 42.890 59.440 43.290 59.840 ;
        RECT 44.890 59.440 45.290 59.840 ;
        RECT 46.890 59.440 47.290 59.840 ;
        RECT 48.890 59.440 49.290 59.840 ;
        RECT 50.890 59.440 51.290 59.840 ;
        RECT 52.890 59.440 53.290 59.840 ;
        RECT 54.890 59.440 55.290 59.840 ;
        RECT 56.890 59.440 57.290 59.840 ;
        RECT 58.890 59.440 59.290 59.840 ;
        RECT 60.890 59.440 61.290 59.840 ;
        RECT 62.890 59.440 63.290 59.840 ;
        RECT 64.890 59.440 65.290 59.840 ;
        RECT 66.890 59.440 67.290 59.840 ;
        RECT 68.890 59.440 69.290 59.840 ;
        RECT 70.890 59.440 71.290 59.840 ;
        RECT 72.890 59.440 73.290 59.840 ;
        RECT 87.825 59.440 88.225 59.840 ;
        RECT 89.825 59.440 90.225 59.840 ;
        RECT 91.825 59.440 92.225 59.840 ;
        RECT 93.825 59.440 94.225 59.840 ;
        RECT 95.825 59.440 96.225 59.840 ;
        RECT 97.825 59.440 98.225 59.840 ;
        RECT 99.825 59.440 100.225 59.840 ;
        RECT 101.825 59.440 102.225 59.840 ;
        RECT 103.825 59.440 104.225 59.840 ;
        RECT 105.825 59.440 106.225 59.840 ;
        RECT 107.825 59.440 108.225 59.840 ;
        RECT 109.825 59.440 110.225 59.840 ;
        RECT 111.825 59.440 112.225 59.840 ;
        RECT 113.825 59.440 114.225 59.840 ;
        RECT 115.825 59.440 116.225 59.840 ;
        RECT 117.825 59.440 118.225 59.840 ;
        RECT 119.825 59.440 120.225 59.840 ;
        RECT 121.825 59.440 122.225 59.840 ;
        RECT 123.825 59.440 124.225 59.840 ;
        RECT 125.825 59.440 126.225 59.840 ;
        RECT 127.825 59.440 128.225 59.840 ;
        RECT 129.825 59.440 130.225 59.840 ;
        RECT 131.825 59.440 132.225 59.840 ;
        RECT 133.825 59.440 134.225 59.840 ;
        RECT 135.825 59.440 136.225 59.840 ;
        RECT 137.825 59.440 138.225 59.840 ;
        RECT 139.825 59.440 140.225 59.840 ;
        RECT 141.825 59.440 142.225 59.840 ;
        RECT 143.825 59.440 144.225 59.840 ;
        RECT 145.825 59.440 146.225 59.840 ;
        RECT 147.825 59.440 148.225 59.840 ;
        RECT 149.825 59.440 150.225 59.840 ;
        RECT 151.825 59.440 152.225 59.840 ;
        RECT 153.825 59.440 154.225 59.840 ;
        RECT 6.890 59.240 8.540 59.440 ;
        RECT 8.890 59.240 22.540 59.440 ;
        RECT 22.890 59.240 38.540 59.440 ;
        RECT 38.890 59.240 46.540 59.440 ;
        RECT 46.890 59.240 50.540 59.440 ;
        RECT 50.890 59.240 52.540 59.440 ;
        RECT 52.890 59.240 54.540 59.440 ;
        RECT 54.890 59.240 60.540 59.440 ;
        RECT 60.890 59.240 64.540 59.440 ;
        RECT 64.890 59.240 74.540 59.440 ;
        RECT 86.575 59.240 96.225 59.440 ;
        RECT 96.575 59.240 100.225 59.440 ;
        RECT 100.575 59.240 106.225 59.440 ;
        RECT 106.575 59.240 108.225 59.440 ;
        RECT 108.575 59.240 110.225 59.440 ;
        RECT 110.575 59.240 114.225 59.440 ;
        RECT 114.575 59.240 122.225 59.440 ;
        RECT 122.575 59.240 138.225 59.440 ;
        RECT 138.575 59.240 152.225 59.440 ;
        RECT 152.575 59.240 154.225 59.440 ;
        RECT 6.890 58.840 7.290 59.240 ;
        RECT 8.890 58.840 9.290 59.240 ;
        RECT 10.890 58.840 11.290 59.240 ;
        RECT 12.890 58.840 13.290 59.240 ;
        RECT 14.890 58.840 15.290 59.240 ;
        RECT 16.890 58.840 17.290 59.240 ;
        RECT 18.890 58.840 19.290 59.240 ;
        RECT 20.890 58.840 21.290 59.240 ;
        RECT 22.890 58.840 23.290 59.240 ;
        RECT 24.890 58.840 25.290 59.240 ;
        RECT 26.890 58.840 27.290 59.240 ;
        RECT 28.890 58.840 29.290 59.240 ;
        RECT 30.890 58.840 31.290 59.240 ;
        RECT 32.890 58.840 33.290 59.240 ;
        RECT 34.890 58.840 35.290 59.240 ;
        RECT 36.890 58.840 37.290 59.240 ;
        RECT 38.890 58.840 39.290 59.240 ;
        RECT 40.890 58.840 41.290 59.240 ;
        RECT 42.890 58.840 43.290 59.240 ;
        RECT 44.890 58.840 45.290 59.240 ;
        RECT 46.890 58.840 47.290 59.240 ;
        RECT 48.890 58.840 49.290 59.240 ;
        RECT 50.890 58.840 51.290 59.240 ;
        RECT 52.890 58.840 53.290 59.240 ;
        RECT 54.890 58.840 55.290 59.240 ;
        RECT 56.890 58.840 57.290 59.240 ;
        RECT 58.890 58.840 59.290 59.240 ;
        RECT 60.890 58.840 61.290 59.240 ;
        RECT 62.890 58.840 63.290 59.240 ;
        RECT 64.890 58.840 65.290 59.240 ;
        RECT 66.890 58.840 67.290 59.240 ;
        RECT 68.890 58.840 69.290 59.240 ;
        RECT 70.890 58.840 71.290 59.240 ;
        RECT 72.890 58.840 73.290 59.240 ;
        RECT 87.825 58.840 88.225 59.240 ;
        RECT 89.825 58.840 90.225 59.240 ;
        RECT 91.825 58.840 92.225 59.240 ;
        RECT 93.825 58.840 94.225 59.240 ;
        RECT 95.825 58.840 96.225 59.240 ;
        RECT 97.825 58.840 98.225 59.240 ;
        RECT 99.825 58.840 100.225 59.240 ;
        RECT 101.825 58.840 102.225 59.240 ;
        RECT 103.825 58.840 104.225 59.240 ;
        RECT 105.825 58.840 106.225 59.240 ;
        RECT 107.825 58.840 108.225 59.240 ;
        RECT 109.825 58.840 110.225 59.240 ;
        RECT 111.825 58.840 112.225 59.240 ;
        RECT 113.825 58.840 114.225 59.240 ;
        RECT 115.825 58.840 116.225 59.240 ;
        RECT 117.825 58.840 118.225 59.240 ;
        RECT 119.825 58.840 120.225 59.240 ;
        RECT 121.825 58.840 122.225 59.240 ;
        RECT 123.825 58.840 124.225 59.240 ;
        RECT 125.825 58.840 126.225 59.240 ;
        RECT 127.825 58.840 128.225 59.240 ;
        RECT 129.825 58.840 130.225 59.240 ;
        RECT 131.825 58.840 132.225 59.240 ;
        RECT 133.825 58.840 134.225 59.240 ;
        RECT 135.825 58.840 136.225 59.240 ;
        RECT 137.825 58.840 138.225 59.240 ;
        RECT 139.825 58.840 140.225 59.240 ;
        RECT 141.825 58.840 142.225 59.240 ;
        RECT 143.825 58.840 144.225 59.240 ;
        RECT 145.825 58.840 146.225 59.240 ;
        RECT 147.825 58.840 148.225 59.240 ;
        RECT 149.825 58.840 150.225 59.240 ;
        RECT 151.825 58.840 152.225 59.240 ;
        RECT 153.825 58.840 154.225 59.240 ;
        RECT 6.960 57.990 7.220 58.840 ;
        RECT 8.990 57.990 9.190 58.840 ;
        RECT 10.990 57.990 11.190 58.840 ;
        RECT 12.990 57.990 13.190 58.840 ;
        RECT 14.990 57.990 15.190 58.840 ;
        RECT 16.990 57.990 17.190 58.840 ;
        RECT 18.990 57.990 19.190 58.840 ;
        RECT 20.990 57.990 21.190 58.840 ;
        RECT 22.990 57.990 23.190 58.840 ;
        RECT 24.990 57.990 25.190 58.840 ;
        RECT 26.990 57.990 27.190 58.840 ;
        RECT 28.990 57.990 29.190 58.840 ;
        RECT 30.990 57.990 31.190 58.840 ;
        RECT 32.990 57.990 33.190 58.840 ;
        RECT 34.990 57.990 35.190 58.840 ;
        RECT 36.990 57.990 37.190 58.840 ;
        RECT 38.990 57.990 39.190 58.840 ;
        RECT 40.990 57.990 41.190 58.840 ;
        RECT 42.990 57.990 43.190 58.840 ;
        RECT 44.990 57.990 45.190 58.840 ;
        RECT 46.990 57.990 47.190 58.840 ;
        RECT 48.990 57.990 49.190 58.840 ;
        RECT 50.990 57.990 51.190 58.840 ;
        RECT 52.990 57.990 53.190 58.840 ;
        RECT 54.990 57.990 55.190 58.840 ;
        RECT 56.990 57.990 57.190 58.840 ;
        RECT 58.990 57.990 59.190 58.840 ;
        RECT 60.990 57.990 61.190 58.840 ;
        RECT 62.990 57.990 63.190 58.840 ;
        RECT 97.925 57.990 98.125 58.840 ;
        RECT 99.925 57.990 100.125 58.840 ;
        RECT 101.925 57.990 102.125 58.840 ;
        RECT 103.925 57.990 104.125 58.840 ;
        RECT 105.925 57.990 106.125 58.840 ;
        RECT 107.925 57.990 108.125 58.840 ;
        RECT 109.925 57.990 110.125 58.840 ;
        RECT 111.925 57.990 112.125 58.840 ;
        RECT 113.925 57.990 114.125 58.840 ;
        RECT 115.925 57.990 116.125 58.840 ;
        RECT 117.925 57.990 118.125 58.840 ;
        RECT 119.925 57.990 120.125 58.840 ;
        RECT 121.925 57.990 122.125 58.840 ;
        RECT 123.925 57.990 124.125 58.840 ;
        RECT 125.925 57.990 126.125 58.840 ;
        RECT 127.925 57.990 128.125 58.840 ;
        RECT 129.925 57.990 130.125 58.840 ;
        RECT 131.925 57.990 132.125 58.840 ;
        RECT 133.925 57.990 134.125 58.840 ;
        RECT 135.925 57.990 136.125 58.840 ;
        RECT 137.925 57.990 138.125 58.840 ;
        RECT 139.925 57.990 140.125 58.840 ;
        RECT 141.925 57.990 142.125 58.840 ;
        RECT 143.925 57.990 144.125 58.840 ;
        RECT 145.925 57.990 146.125 58.840 ;
        RECT 147.925 57.990 148.125 58.840 ;
        RECT 149.925 57.990 150.125 58.840 ;
        RECT 151.925 57.990 152.125 58.840 ;
        RECT 153.895 57.990 154.155 58.840 ;
        RECT 6.890 57.590 7.290 57.990 ;
        RECT 8.890 57.590 9.290 57.990 ;
        RECT 10.890 57.590 11.290 57.990 ;
        RECT 12.890 57.590 13.290 57.990 ;
        RECT 14.890 57.590 15.290 57.990 ;
        RECT 16.890 57.590 17.290 57.990 ;
        RECT 18.890 57.590 19.290 57.990 ;
        RECT 20.890 57.590 21.290 57.990 ;
        RECT 22.890 57.590 23.290 57.990 ;
        RECT 24.890 57.590 25.290 57.990 ;
        RECT 26.890 57.590 27.290 57.990 ;
        RECT 28.890 57.590 29.290 57.990 ;
        RECT 30.890 57.590 31.290 57.990 ;
        RECT 32.890 57.590 33.290 57.990 ;
        RECT 34.890 57.590 35.290 57.990 ;
        RECT 36.890 57.590 37.290 57.990 ;
        RECT 38.890 57.590 39.290 57.990 ;
        RECT 40.890 57.590 41.290 57.990 ;
        RECT 42.890 57.590 43.290 57.990 ;
        RECT 44.890 57.590 45.290 57.990 ;
        RECT 46.890 57.590 47.290 57.990 ;
        RECT 48.890 57.590 49.290 57.990 ;
        RECT 50.890 57.590 51.290 57.990 ;
        RECT 52.890 57.590 53.290 57.990 ;
        RECT 54.890 57.590 55.290 57.990 ;
        RECT 56.890 57.590 57.290 57.990 ;
        RECT 58.890 57.590 59.290 57.990 ;
        RECT 60.890 57.590 61.290 57.990 ;
        RECT 62.890 57.590 63.290 57.990 ;
        RECT 64.890 57.590 65.290 57.990 ;
        RECT 66.890 57.590 67.290 57.990 ;
        RECT 68.890 57.590 69.290 57.990 ;
        RECT 70.890 57.590 71.290 57.990 ;
        RECT 72.890 57.590 73.290 57.990 ;
        RECT 77.180 57.590 77.600 57.670 ;
        RECT 6.890 57.390 8.540 57.590 ;
        RECT 8.890 57.390 22.540 57.590 ;
        RECT 22.890 57.390 38.540 57.590 ;
        RECT 38.890 57.390 46.540 57.590 ;
        RECT 46.890 57.390 50.540 57.590 ;
        RECT 50.890 57.390 52.540 57.590 ;
        RECT 52.890 57.390 54.540 57.590 ;
        RECT 54.890 57.390 60.540 57.590 ;
        RECT 60.890 57.390 77.600 57.590 ;
        RECT 6.890 56.990 7.290 57.390 ;
        RECT 8.890 56.990 9.290 57.390 ;
        RECT 10.890 56.990 11.290 57.390 ;
        RECT 12.890 56.990 13.290 57.390 ;
        RECT 14.890 56.990 15.290 57.390 ;
        RECT 16.890 56.990 17.290 57.390 ;
        RECT 18.890 56.990 19.290 57.390 ;
        RECT 20.890 56.990 21.290 57.390 ;
        RECT 22.890 56.990 23.290 57.390 ;
        RECT 24.890 56.990 25.290 57.390 ;
        RECT 26.890 56.990 27.290 57.390 ;
        RECT 28.890 56.990 29.290 57.390 ;
        RECT 30.890 56.990 31.290 57.390 ;
        RECT 32.890 56.990 33.290 57.390 ;
        RECT 34.890 56.990 35.290 57.390 ;
        RECT 36.890 56.990 37.290 57.390 ;
        RECT 38.890 56.990 39.290 57.390 ;
        RECT 40.890 56.990 41.290 57.390 ;
        RECT 42.890 56.990 43.290 57.390 ;
        RECT 44.890 56.990 45.290 57.390 ;
        RECT 46.890 56.990 47.290 57.390 ;
        RECT 48.890 56.990 49.290 57.390 ;
        RECT 50.890 56.990 51.290 57.390 ;
        RECT 52.890 56.990 53.290 57.390 ;
        RECT 54.890 56.990 55.290 57.390 ;
        RECT 56.890 56.990 57.290 57.390 ;
        RECT 58.890 56.990 59.290 57.390 ;
        RECT 60.890 56.990 61.290 57.390 ;
        RECT 62.890 56.990 63.290 57.390 ;
        RECT 64.890 56.990 65.290 57.390 ;
        RECT 66.890 56.990 67.290 57.390 ;
        RECT 68.890 56.990 69.290 57.390 ;
        RECT 70.890 56.990 71.290 57.390 ;
        RECT 72.890 56.990 73.290 57.390 ;
        RECT 77.180 57.310 77.600 57.390 ;
        RECT 83.515 57.590 83.935 57.670 ;
        RECT 87.825 57.590 88.225 57.990 ;
        RECT 89.825 57.590 90.225 57.990 ;
        RECT 91.825 57.590 92.225 57.990 ;
        RECT 93.825 57.590 94.225 57.990 ;
        RECT 95.825 57.590 96.225 57.990 ;
        RECT 97.825 57.590 98.225 57.990 ;
        RECT 99.825 57.590 100.225 57.990 ;
        RECT 101.825 57.590 102.225 57.990 ;
        RECT 103.825 57.590 104.225 57.990 ;
        RECT 105.825 57.590 106.225 57.990 ;
        RECT 107.825 57.590 108.225 57.990 ;
        RECT 109.825 57.590 110.225 57.990 ;
        RECT 111.825 57.590 112.225 57.990 ;
        RECT 113.825 57.590 114.225 57.990 ;
        RECT 115.825 57.590 116.225 57.990 ;
        RECT 117.825 57.590 118.225 57.990 ;
        RECT 119.825 57.590 120.225 57.990 ;
        RECT 121.825 57.590 122.225 57.990 ;
        RECT 123.825 57.590 124.225 57.990 ;
        RECT 125.825 57.590 126.225 57.990 ;
        RECT 127.825 57.590 128.225 57.990 ;
        RECT 129.825 57.590 130.225 57.990 ;
        RECT 131.825 57.590 132.225 57.990 ;
        RECT 133.825 57.590 134.225 57.990 ;
        RECT 135.825 57.590 136.225 57.990 ;
        RECT 137.825 57.590 138.225 57.990 ;
        RECT 139.825 57.590 140.225 57.990 ;
        RECT 141.825 57.590 142.225 57.990 ;
        RECT 143.825 57.590 144.225 57.990 ;
        RECT 145.825 57.590 146.225 57.990 ;
        RECT 147.825 57.590 148.225 57.990 ;
        RECT 149.825 57.590 150.225 57.990 ;
        RECT 151.825 57.590 152.225 57.990 ;
        RECT 153.825 57.590 154.225 57.990 ;
        RECT 83.515 57.390 100.225 57.590 ;
        RECT 100.575 57.390 106.225 57.590 ;
        RECT 106.575 57.390 108.225 57.590 ;
        RECT 108.575 57.390 110.225 57.590 ;
        RECT 110.575 57.390 114.225 57.590 ;
        RECT 114.575 57.390 122.225 57.590 ;
        RECT 122.575 57.390 138.225 57.590 ;
        RECT 138.575 57.390 152.225 57.590 ;
        RECT 152.575 57.390 154.225 57.590 ;
        RECT 83.515 57.310 83.935 57.390 ;
        RECT 87.825 56.990 88.225 57.390 ;
        RECT 89.825 56.990 90.225 57.390 ;
        RECT 91.825 56.990 92.225 57.390 ;
        RECT 93.825 56.990 94.225 57.390 ;
        RECT 95.825 56.990 96.225 57.390 ;
        RECT 97.825 56.990 98.225 57.390 ;
        RECT 99.825 56.990 100.225 57.390 ;
        RECT 101.825 56.990 102.225 57.390 ;
        RECT 103.825 56.990 104.225 57.390 ;
        RECT 105.825 56.990 106.225 57.390 ;
        RECT 107.825 56.990 108.225 57.390 ;
        RECT 109.825 56.990 110.225 57.390 ;
        RECT 111.825 56.990 112.225 57.390 ;
        RECT 113.825 56.990 114.225 57.390 ;
        RECT 115.825 56.990 116.225 57.390 ;
        RECT 117.825 56.990 118.225 57.390 ;
        RECT 119.825 56.990 120.225 57.390 ;
        RECT 121.825 56.990 122.225 57.390 ;
        RECT 123.825 56.990 124.225 57.390 ;
        RECT 125.825 56.990 126.225 57.390 ;
        RECT 127.825 56.990 128.225 57.390 ;
        RECT 129.825 56.990 130.225 57.390 ;
        RECT 131.825 56.990 132.225 57.390 ;
        RECT 133.825 56.990 134.225 57.390 ;
        RECT 135.825 56.990 136.225 57.390 ;
        RECT 137.825 56.990 138.225 57.390 ;
        RECT 139.825 56.990 140.225 57.390 ;
        RECT 141.825 56.990 142.225 57.390 ;
        RECT 143.825 56.990 144.225 57.390 ;
        RECT 145.825 56.990 146.225 57.390 ;
        RECT 147.825 56.990 148.225 57.390 ;
        RECT 149.825 56.990 150.225 57.390 ;
        RECT 151.825 56.990 152.225 57.390 ;
        RECT 153.825 56.990 154.225 57.390 ;
        RECT 6.960 56.140 7.220 56.990 ;
        RECT 8.990 56.140 9.190 56.990 ;
        RECT 10.990 56.140 11.190 56.990 ;
        RECT 12.990 56.140 13.190 56.990 ;
        RECT 14.990 56.140 15.190 56.990 ;
        RECT 16.990 56.140 17.190 56.990 ;
        RECT 18.990 56.140 19.190 56.990 ;
        RECT 20.990 56.140 21.190 56.990 ;
        RECT 22.990 56.140 23.190 56.990 ;
        RECT 24.990 56.140 25.190 56.990 ;
        RECT 26.990 56.140 27.190 56.990 ;
        RECT 28.990 56.140 29.190 56.990 ;
        RECT 30.990 56.140 31.190 56.990 ;
        RECT 32.990 56.140 33.190 56.990 ;
        RECT 34.990 56.140 35.190 56.990 ;
        RECT 36.990 56.140 37.190 56.990 ;
        RECT 38.990 56.140 39.190 56.990 ;
        RECT 40.990 56.140 41.190 56.990 ;
        RECT 42.990 56.140 43.190 56.990 ;
        RECT 44.990 56.140 45.190 56.990 ;
        RECT 46.990 56.140 47.190 56.990 ;
        RECT 48.990 56.140 49.190 56.990 ;
        RECT 50.990 56.140 51.190 56.990 ;
        RECT 52.990 56.140 53.190 56.990 ;
        RECT 54.990 56.140 55.190 56.990 ;
        RECT 56.990 56.140 57.190 56.990 ;
        RECT 58.990 56.140 59.190 56.990 ;
        RECT 101.925 56.140 102.125 56.990 ;
        RECT 103.925 56.140 104.125 56.990 ;
        RECT 105.925 56.140 106.125 56.990 ;
        RECT 107.925 56.140 108.125 56.990 ;
        RECT 109.925 56.140 110.125 56.990 ;
        RECT 111.925 56.140 112.125 56.990 ;
        RECT 113.925 56.140 114.125 56.990 ;
        RECT 115.925 56.140 116.125 56.990 ;
        RECT 117.925 56.140 118.125 56.990 ;
        RECT 119.925 56.140 120.125 56.990 ;
        RECT 121.925 56.140 122.125 56.990 ;
        RECT 123.925 56.140 124.125 56.990 ;
        RECT 125.925 56.140 126.125 56.990 ;
        RECT 127.925 56.140 128.125 56.990 ;
        RECT 129.925 56.140 130.125 56.990 ;
        RECT 131.925 56.140 132.125 56.990 ;
        RECT 133.925 56.140 134.125 56.990 ;
        RECT 135.925 56.140 136.125 56.990 ;
        RECT 137.925 56.140 138.125 56.990 ;
        RECT 139.925 56.140 140.125 56.990 ;
        RECT 141.925 56.140 142.125 56.990 ;
        RECT 143.925 56.140 144.125 56.990 ;
        RECT 145.925 56.140 146.125 56.990 ;
        RECT 147.925 56.140 148.125 56.990 ;
        RECT 149.925 56.140 150.125 56.990 ;
        RECT 151.925 56.140 152.125 56.990 ;
        RECT 153.895 56.140 154.155 56.990 ;
        RECT 6.890 55.740 7.290 56.140 ;
        RECT 8.890 55.740 9.290 56.140 ;
        RECT 10.890 55.740 11.290 56.140 ;
        RECT 12.890 55.740 13.290 56.140 ;
        RECT 14.890 55.740 15.290 56.140 ;
        RECT 16.890 55.740 17.290 56.140 ;
        RECT 18.890 55.740 19.290 56.140 ;
        RECT 20.890 55.740 21.290 56.140 ;
        RECT 22.890 55.740 23.290 56.140 ;
        RECT 24.890 55.740 25.290 56.140 ;
        RECT 26.890 55.740 27.290 56.140 ;
        RECT 28.890 55.740 29.290 56.140 ;
        RECT 30.890 55.740 31.290 56.140 ;
        RECT 32.890 55.740 33.290 56.140 ;
        RECT 34.890 55.740 35.290 56.140 ;
        RECT 36.890 55.740 37.290 56.140 ;
        RECT 38.890 55.740 39.290 56.140 ;
        RECT 40.890 55.740 41.290 56.140 ;
        RECT 42.890 55.740 43.290 56.140 ;
        RECT 44.890 55.740 45.290 56.140 ;
        RECT 46.890 55.740 47.290 56.140 ;
        RECT 48.890 55.740 49.290 56.140 ;
        RECT 50.890 55.740 51.290 56.140 ;
        RECT 52.890 55.740 53.290 56.140 ;
        RECT 54.890 55.740 55.290 56.140 ;
        RECT 56.890 55.740 57.290 56.140 ;
        RECT 58.890 55.740 59.290 56.140 ;
        RECT 60.890 55.740 61.290 56.140 ;
        RECT 62.890 55.740 63.290 56.140 ;
        RECT 64.890 55.740 65.290 56.140 ;
        RECT 66.890 55.740 67.290 56.140 ;
        RECT 68.890 55.740 69.290 56.140 ;
        RECT 70.890 55.740 71.290 56.140 ;
        RECT 72.890 55.740 73.290 56.140 ;
        RECT 76.730 55.740 77.150 55.820 ;
        RECT 6.890 55.540 8.540 55.740 ;
        RECT 8.890 55.540 22.540 55.740 ;
        RECT 22.890 55.540 38.540 55.740 ;
        RECT 38.890 55.540 46.540 55.740 ;
        RECT 46.890 55.540 50.540 55.740 ;
        RECT 50.890 55.540 52.540 55.740 ;
        RECT 52.890 55.540 54.540 55.740 ;
        RECT 54.890 55.540 77.150 55.740 ;
        RECT 6.890 55.140 7.290 55.540 ;
        RECT 8.890 55.140 9.290 55.540 ;
        RECT 10.890 55.140 11.290 55.540 ;
        RECT 12.890 55.140 13.290 55.540 ;
        RECT 14.890 55.140 15.290 55.540 ;
        RECT 16.890 55.140 17.290 55.540 ;
        RECT 18.890 55.140 19.290 55.540 ;
        RECT 20.890 55.140 21.290 55.540 ;
        RECT 22.890 55.140 23.290 55.540 ;
        RECT 24.890 55.140 25.290 55.540 ;
        RECT 26.890 55.140 27.290 55.540 ;
        RECT 28.890 55.140 29.290 55.540 ;
        RECT 30.890 55.140 31.290 55.540 ;
        RECT 32.890 55.140 33.290 55.540 ;
        RECT 34.890 55.140 35.290 55.540 ;
        RECT 36.890 55.140 37.290 55.540 ;
        RECT 38.890 55.140 39.290 55.540 ;
        RECT 40.890 55.140 41.290 55.540 ;
        RECT 42.890 55.140 43.290 55.540 ;
        RECT 44.890 55.140 45.290 55.540 ;
        RECT 46.890 55.140 47.290 55.540 ;
        RECT 48.890 55.140 49.290 55.540 ;
        RECT 50.890 55.140 51.290 55.540 ;
        RECT 52.890 55.140 53.290 55.540 ;
        RECT 54.890 55.140 55.290 55.540 ;
        RECT 56.890 55.140 57.290 55.540 ;
        RECT 58.890 55.140 59.290 55.540 ;
        RECT 60.890 55.140 61.290 55.540 ;
        RECT 62.890 55.140 63.290 55.540 ;
        RECT 64.890 55.140 65.290 55.540 ;
        RECT 66.890 55.140 67.290 55.540 ;
        RECT 68.890 55.140 69.290 55.540 ;
        RECT 70.890 55.140 71.290 55.540 ;
        RECT 72.890 55.140 73.290 55.540 ;
        RECT 76.730 55.460 77.150 55.540 ;
        RECT 83.965 55.740 84.385 55.820 ;
        RECT 87.825 55.740 88.225 56.140 ;
        RECT 89.825 55.740 90.225 56.140 ;
        RECT 91.825 55.740 92.225 56.140 ;
        RECT 93.825 55.740 94.225 56.140 ;
        RECT 95.825 55.740 96.225 56.140 ;
        RECT 97.825 55.740 98.225 56.140 ;
        RECT 99.825 55.740 100.225 56.140 ;
        RECT 101.825 55.740 102.225 56.140 ;
        RECT 103.825 55.740 104.225 56.140 ;
        RECT 105.825 55.740 106.225 56.140 ;
        RECT 107.825 55.740 108.225 56.140 ;
        RECT 109.825 55.740 110.225 56.140 ;
        RECT 111.825 55.740 112.225 56.140 ;
        RECT 113.825 55.740 114.225 56.140 ;
        RECT 115.825 55.740 116.225 56.140 ;
        RECT 117.825 55.740 118.225 56.140 ;
        RECT 119.825 55.740 120.225 56.140 ;
        RECT 121.825 55.740 122.225 56.140 ;
        RECT 123.825 55.740 124.225 56.140 ;
        RECT 125.825 55.740 126.225 56.140 ;
        RECT 127.825 55.740 128.225 56.140 ;
        RECT 129.825 55.740 130.225 56.140 ;
        RECT 131.825 55.740 132.225 56.140 ;
        RECT 133.825 55.740 134.225 56.140 ;
        RECT 135.825 55.740 136.225 56.140 ;
        RECT 137.825 55.740 138.225 56.140 ;
        RECT 139.825 55.740 140.225 56.140 ;
        RECT 141.825 55.740 142.225 56.140 ;
        RECT 143.825 55.740 144.225 56.140 ;
        RECT 145.825 55.740 146.225 56.140 ;
        RECT 147.825 55.740 148.225 56.140 ;
        RECT 149.825 55.740 150.225 56.140 ;
        RECT 151.825 55.740 152.225 56.140 ;
        RECT 153.825 55.740 154.225 56.140 ;
        RECT 83.965 55.540 106.225 55.740 ;
        RECT 106.575 55.540 108.225 55.740 ;
        RECT 108.575 55.540 110.225 55.740 ;
        RECT 110.575 55.540 114.225 55.740 ;
        RECT 114.575 55.540 122.225 55.740 ;
        RECT 122.575 55.540 138.225 55.740 ;
        RECT 138.575 55.540 152.225 55.740 ;
        RECT 152.575 55.540 154.225 55.740 ;
        RECT 83.965 55.460 84.385 55.540 ;
        RECT 87.825 55.140 88.225 55.540 ;
        RECT 89.825 55.140 90.225 55.540 ;
        RECT 91.825 55.140 92.225 55.540 ;
        RECT 93.825 55.140 94.225 55.540 ;
        RECT 95.825 55.140 96.225 55.540 ;
        RECT 97.825 55.140 98.225 55.540 ;
        RECT 99.825 55.140 100.225 55.540 ;
        RECT 101.825 55.140 102.225 55.540 ;
        RECT 103.825 55.140 104.225 55.540 ;
        RECT 105.825 55.140 106.225 55.540 ;
        RECT 107.825 55.140 108.225 55.540 ;
        RECT 109.825 55.140 110.225 55.540 ;
        RECT 111.825 55.140 112.225 55.540 ;
        RECT 113.825 55.140 114.225 55.540 ;
        RECT 115.825 55.140 116.225 55.540 ;
        RECT 117.825 55.140 118.225 55.540 ;
        RECT 119.825 55.140 120.225 55.540 ;
        RECT 121.825 55.140 122.225 55.540 ;
        RECT 123.825 55.140 124.225 55.540 ;
        RECT 125.825 55.140 126.225 55.540 ;
        RECT 127.825 55.140 128.225 55.540 ;
        RECT 129.825 55.140 130.225 55.540 ;
        RECT 131.825 55.140 132.225 55.540 ;
        RECT 133.825 55.140 134.225 55.540 ;
        RECT 135.825 55.140 136.225 55.540 ;
        RECT 137.825 55.140 138.225 55.540 ;
        RECT 139.825 55.140 140.225 55.540 ;
        RECT 141.825 55.140 142.225 55.540 ;
        RECT 143.825 55.140 144.225 55.540 ;
        RECT 145.825 55.140 146.225 55.540 ;
        RECT 147.825 55.140 148.225 55.540 ;
        RECT 149.825 55.140 150.225 55.540 ;
        RECT 151.825 55.140 152.225 55.540 ;
        RECT 153.825 55.140 154.225 55.540 ;
        RECT 6.960 54.290 7.220 55.140 ;
        RECT 8.990 54.290 9.190 55.140 ;
        RECT 10.990 54.290 11.190 55.140 ;
        RECT 12.990 54.290 13.190 55.140 ;
        RECT 14.990 54.290 15.190 55.140 ;
        RECT 16.990 54.290 17.190 55.140 ;
        RECT 18.990 54.290 19.190 55.140 ;
        RECT 20.990 54.290 21.190 55.140 ;
        RECT 22.990 54.290 23.190 55.140 ;
        RECT 24.990 54.290 25.190 55.140 ;
        RECT 26.990 54.290 27.190 55.140 ;
        RECT 28.990 54.290 29.190 55.140 ;
        RECT 30.990 54.290 31.190 55.140 ;
        RECT 32.990 54.290 33.190 55.140 ;
        RECT 34.990 54.290 35.190 55.140 ;
        RECT 36.990 54.290 37.190 55.140 ;
        RECT 38.990 54.290 39.190 55.140 ;
        RECT 40.990 54.290 41.190 55.140 ;
        RECT 42.990 54.290 43.190 55.140 ;
        RECT 44.990 54.290 45.190 55.140 ;
        RECT 46.990 54.290 47.190 55.140 ;
        RECT 48.990 54.290 49.190 55.140 ;
        RECT 50.990 54.290 51.190 55.140 ;
        RECT 52.990 54.290 53.190 55.140 ;
        RECT 54.990 54.290 55.190 55.140 ;
        RECT 56.990 54.290 57.190 55.140 ;
        RECT 58.990 54.290 59.190 55.140 ;
        RECT 60.990 54.290 61.190 55.140 ;
        RECT 62.990 54.290 63.190 55.140 ;
        RECT 64.990 54.290 65.190 55.140 ;
        RECT 66.990 54.290 67.190 55.140 ;
        RECT 68.990 54.290 69.190 55.140 ;
        RECT 70.990 54.290 71.190 55.140 ;
        RECT 89.925 54.290 90.125 55.140 ;
        RECT 91.925 54.290 92.125 55.140 ;
        RECT 93.925 54.290 94.125 55.140 ;
        RECT 95.925 54.290 96.125 55.140 ;
        RECT 97.925 54.290 98.125 55.140 ;
        RECT 99.925 54.290 100.125 55.140 ;
        RECT 101.925 54.290 102.125 55.140 ;
        RECT 103.925 54.290 104.125 55.140 ;
        RECT 105.925 54.290 106.125 55.140 ;
        RECT 107.925 54.290 108.125 55.140 ;
        RECT 109.925 54.290 110.125 55.140 ;
        RECT 111.925 54.290 112.125 55.140 ;
        RECT 113.925 54.290 114.125 55.140 ;
        RECT 115.925 54.290 116.125 55.140 ;
        RECT 117.925 54.290 118.125 55.140 ;
        RECT 119.925 54.290 120.125 55.140 ;
        RECT 121.925 54.290 122.125 55.140 ;
        RECT 123.925 54.290 124.125 55.140 ;
        RECT 125.925 54.290 126.125 55.140 ;
        RECT 127.925 54.290 128.125 55.140 ;
        RECT 129.925 54.290 130.125 55.140 ;
        RECT 131.925 54.290 132.125 55.140 ;
        RECT 133.925 54.290 134.125 55.140 ;
        RECT 135.925 54.290 136.125 55.140 ;
        RECT 137.925 54.290 138.125 55.140 ;
        RECT 139.925 54.290 140.125 55.140 ;
        RECT 141.925 54.290 142.125 55.140 ;
        RECT 143.925 54.290 144.125 55.140 ;
        RECT 145.925 54.290 146.125 55.140 ;
        RECT 147.925 54.290 148.125 55.140 ;
        RECT 149.925 54.290 150.125 55.140 ;
        RECT 151.925 54.290 152.125 55.140 ;
        RECT 153.895 54.290 154.155 55.140 ;
        RECT 6.890 53.890 7.290 54.290 ;
        RECT 8.890 53.890 9.290 54.290 ;
        RECT 10.890 53.890 11.290 54.290 ;
        RECT 12.890 53.890 13.290 54.290 ;
        RECT 14.890 53.890 15.290 54.290 ;
        RECT 16.890 53.890 17.290 54.290 ;
        RECT 18.890 53.890 19.290 54.290 ;
        RECT 20.890 53.890 21.290 54.290 ;
        RECT 22.890 53.890 23.290 54.290 ;
        RECT 24.890 53.890 25.290 54.290 ;
        RECT 26.890 53.890 27.290 54.290 ;
        RECT 28.890 53.890 29.290 54.290 ;
        RECT 30.890 53.890 31.290 54.290 ;
        RECT 32.890 53.890 33.290 54.290 ;
        RECT 34.890 53.890 35.290 54.290 ;
        RECT 36.890 53.890 37.290 54.290 ;
        RECT 38.890 53.890 39.290 54.290 ;
        RECT 40.890 53.890 41.290 54.290 ;
        RECT 42.890 53.890 43.290 54.290 ;
        RECT 44.890 53.890 45.290 54.290 ;
        RECT 46.890 53.890 47.290 54.290 ;
        RECT 48.890 53.890 49.290 54.290 ;
        RECT 50.890 53.890 51.290 54.290 ;
        RECT 52.890 53.890 53.290 54.290 ;
        RECT 54.890 53.890 55.290 54.290 ;
        RECT 56.890 53.890 57.290 54.290 ;
        RECT 58.890 53.890 59.290 54.290 ;
        RECT 60.890 53.890 61.290 54.290 ;
        RECT 62.890 53.890 63.290 54.290 ;
        RECT 64.890 53.890 65.290 54.290 ;
        RECT 66.890 53.890 67.290 54.290 ;
        RECT 68.890 53.890 69.290 54.290 ;
        RECT 70.890 53.890 71.290 54.290 ;
        RECT 72.890 53.890 73.290 54.290 ;
        RECT 87.825 53.890 88.225 54.290 ;
        RECT 89.825 53.890 90.225 54.290 ;
        RECT 91.825 53.890 92.225 54.290 ;
        RECT 93.825 53.890 94.225 54.290 ;
        RECT 95.825 53.890 96.225 54.290 ;
        RECT 97.825 53.890 98.225 54.290 ;
        RECT 99.825 53.890 100.225 54.290 ;
        RECT 101.825 53.890 102.225 54.290 ;
        RECT 103.825 53.890 104.225 54.290 ;
        RECT 105.825 53.890 106.225 54.290 ;
        RECT 107.825 53.890 108.225 54.290 ;
        RECT 109.825 53.890 110.225 54.290 ;
        RECT 111.825 53.890 112.225 54.290 ;
        RECT 113.825 53.890 114.225 54.290 ;
        RECT 115.825 53.890 116.225 54.290 ;
        RECT 117.825 53.890 118.225 54.290 ;
        RECT 119.825 53.890 120.225 54.290 ;
        RECT 121.825 53.890 122.225 54.290 ;
        RECT 123.825 53.890 124.225 54.290 ;
        RECT 125.825 53.890 126.225 54.290 ;
        RECT 127.825 53.890 128.225 54.290 ;
        RECT 129.825 53.890 130.225 54.290 ;
        RECT 131.825 53.890 132.225 54.290 ;
        RECT 133.825 53.890 134.225 54.290 ;
        RECT 135.825 53.890 136.225 54.290 ;
        RECT 137.825 53.890 138.225 54.290 ;
        RECT 139.825 53.890 140.225 54.290 ;
        RECT 141.825 53.890 142.225 54.290 ;
        RECT 143.825 53.890 144.225 54.290 ;
        RECT 145.825 53.890 146.225 54.290 ;
        RECT 147.825 53.890 148.225 54.290 ;
        RECT 149.825 53.890 150.225 54.290 ;
        RECT 151.825 53.890 152.225 54.290 ;
        RECT 153.825 53.890 154.225 54.290 ;
        RECT 6.890 53.690 8.540 53.890 ;
        RECT 8.890 53.690 22.540 53.890 ;
        RECT 22.890 53.690 38.540 53.890 ;
        RECT 38.890 53.690 46.540 53.890 ;
        RECT 46.890 53.690 50.540 53.890 ;
        RECT 50.890 53.690 52.540 53.890 ;
        RECT 52.890 53.690 54.540 53.890 ;
        RECT 54.890 53.690 74.540 53.890 ;
        RECT 86.575 53.690 106.225 53.890 ;
        RECT 106.575 53.690 108.225 53.890 ;
        RECT 108.575 53.690 110.225 53.890 ;
        RECT 110.575 53.690 114.225 53.890 ;
        RECT 114.575 53.690 122.225 53.890 ;
        RECT 122.575 53.690 138.225 53.890 ;
        RECT 138.575 53.690 152.225 53.890 ;
        RECT 152.575 53.690 154.225 53.890 ;
        RECT 6.890 53.290 7.290 53.690 ;
        RECT 8.890 53.290 9.290 53.690 ;
        RECT 10.890 53.290 11.290 53.690 ;
        RECT 12.890 53.290 13.290 53.690 ;
        RECT 14.890 53.290 15.290 53.690 ;
        RECT 16.890 53.290 17.290 53.690 ;
        RECT 18.890 53.290 19.290 53.690 ;
        RECT 20.890 53.290 21.290 53.690 ;
        RECT 22.890 53.290 23.290 53.690 ;
        RECT 24.890 53.290 25.290 53.690 ;
        RECT 26.890 53.290 27.290 53.690 ;
        RECT 28.890 53.290 29.290 53.690 ;
        RECT 30.890 53.290 31.290 53.690 ;
        RECT 32.890 53.290 33.290 53.690 ;
        RECT 34.890 53.290 35.290 53.690 ;
        RECT 36.890 53.290 37.290 53.690 ;
        RECT 38.890 53.290 39.290 53.690 ;
        RECT 40.890 53.290 41.290 53.690 ;
        RECT 42.890 53.290 43.290 53.690 ;
        RECT 44.890 53.290 45.290 53.690 ;
        RECT 46.890 53.290 47.290 53.690 ;
        RECT 48.890 53.290 49.290 53.690 ;
        RECT 50.890 53.290 51.290 53.690 ;
        RECT 52.890 53.290 53.290 53.690 ;
        RECT 54.890 53.290 55.290 53.690 ;
        RECT 56.890 53.290 57.290 53.690 ;
        RECT 58.890 53.290 59.290 53.690 ;
        RECT 60.890 53.290 61.290 53.690 ;
        RECT 62.890 53.290 63.290 53.690 ;
        RECT 64.890 53.290 65.290 53.690 ;
        RECT 66.890 53.290 67.290 53.690 ;
        RECT 68.890 53.290 69.290 53.690 ;
        RECT 70.890 53.290 71.290 53.690 ;
        RECT 72.890 53.290 73.290 53.690 ;
        RECT 87.825 53.290 88.225 53.690 ;
        RECT 89.825 53.290 90.225 53.690 ;
        RECT 91.825 53.290 92.225 53.690 ;
        RECT 93.825 53.290 94.225 53.690 ;
        RECT 95.825 53.290 96.225 53.690 ;
        RECT 97.825 53.290 98.225 53.690 ;
        RECT 99.825 53.290 100.225 53.690 ;
        RECT 101.825 53.290 102.225 53.690 ;
        RECT 103.825 53.290 104.225 53.690 ;
        RECT 105.825 53.290 106.225 53.690 ;
        RECT 107.825 53.290 108.225 53.690 ;
        RECT 109.825 53.290 110.225 53.690 ;
        RECT 111.825 53.290 112.225 53.690 ;
        RECT 113.825 53.290 114.225 53.690 ;
        RECT 115.825 53.290 116.225 53.690 ;
        RECT 117.825 53.290 118.225 53.690 ;
        RECT 119.825 53.290 120.225 53.690 ;
        RECT 121.825 53.290 122.225 53.690 ;
        RECT 123.825 53.290 124.225 53.690 ;
        RECT 125.825 53.290 126.225 53.690 ;
        RECT 127.825 53.290 128.225 53.690 ;
        RECT 129.825 53.290 130.225 53.690 ;
        RECT 131.825 53.290 132.225 53.690 ;
        RECT 133.825 53.290 134.225 53.690 ;
        RECT 135.825 53.290 136.225 53.690 ;
        RECT 137.825 53.290 138.225 53.690 ;
        RECT 139.825 53.290 140.225 53.690 ;
        RECT 141.825 53.290 142.225 53.690 ;
        RECT 143.825 53.290 144.225 53.690 ;
        RECT 145.825 53.290 146.225 53.690 ;
        RECT 147.825 53.290 148.225 53.690 ;
        RECT 149.825 53.290 150.225 53.690 ;
        RECT 151.825 53.290 152.225 53.690 ;
        RECT 153.825 53.290 154.225 53.690 ;
        RECT 6.960 52.440 7.220 53.290 ;
        RECT 8.990 52.440 9.190 53.290 ;
        RECT 10.990 52.440 11.190 53.290 ;
        RECT 12.990 52.440 13.190 53.290 ;
        RECT 14.990 52.440 15.190 53.290 ;
        RECT 16.990 52.440 17.190 53.290 ;
        RECT 18.990 52.440 19.190 53.290 ;
        RECT 20.990 52.440 21.190 53.290 ;
        RECT 22.990 52.440 23.190 53.290 ;
        RECT 24.990 52.440 25.190 53.290 ;
        RECT 26.990 52.440 27.190 53.290 ;
        RECT 28.990 52.440 29.190 53.290 ;
        RECT 30.990 52.440 31.190 53.290 ;
        RECT 32.990 52.440 33.190 53.290 ;
        RECT 34.990 52.440 35.190 53.290 ;
        RECT 36.990 52.440 37.190 53.290 ;
        RECT 38.990 52.440 39.190 53.290 ;
        RECT 40.990 52.440 41.190 53.290 ;
        RECT 42.990 52.440 43.190 53.290 ;
        RECT 44.990 52.440 45.190 53.290 ;
        RECT 46.990 52.440 47.190 53.290 ;
        RECT 48.990 52.440 49.190 53.290 ;
        RECT 50.990 52.440 51.190 53.290 ;
        RECT 52.990 52.440 53.190 53.290 ;
        RECT 107.925 52.440 108.125 53.290 ;
        RECT 109.925 52.440 110.125 53.290 ;
        RECT 111.925 52.440 112.125 53.290 ;
        RECT 113.925 52.440 114.125 53.290 ;
        RECT 115.925 52.440 116.125 53.290 ;
        RECT 117.925 52.440 118.125 53.290 ;
        RECT 119.925 52.440 120.125 53.290 ;
        RECT 121.925 52.440 122.125 53.290 ;
        RECT 123.925 52.440 124.125 53.290 ;
        RECT 125.925 52.440 126.125 53.290 ;
        RECT 127.925 52.440 128.125 53.290 ;
        RECT 129.925 52.440 130.125 53.290 ;
        RECT 131.925 52.440 132.125 53.290 ;
        RECT 133.925 52.440 134.125 53.290 ;
        RECT 135.925 52.440 136.125 53.290 ;
        RECT 137.925 52.440 138.125 53.290 ;
        RECT 139.925 52.440 140.125 53.290 ;
        RECT 141.925 52.440 142.125 53.290 ;
        RECT 143.925 52.440 144.125 53.290 ;
        RECT 145.925 52.440 146.125 53.290 ;
        RECT 147.925 52.440 148.125 53.290 ;
        RECT 149.925 52.440 150.125 53.290 ;
        RECT 151.925 52.440 152.125 53.290 ;
        RECT 153.895 52.440 154.155 53.290 ;
        RECT 6.890 52.040 7.290 52.440 ;
        RECT 8.890 52.040 9.290 52.440 ;
        RECT 10.890 52.040 11.290 52.440 ;
        RECT 12.890 52.040 13.290 52.440 ;
        RECT 14.890 52.040 15.290 52.440 ;
        RECT 16.890 52.040 17.290 52.440 ;
        RECT 18.890 52.040 19.290 52.440 ;
        RECT 20.890 52.040 21.290 52.440 ;
        RECT 22.890 52.040 23.290 52.440 ;
        RECT 24.890 52.040 25.290 52.440 ;
        RECT 26.890 52.040 27.290 52.440 ;
        RECT 28.890 52.040 29.290 52.440 ;
        RECT 30.890 52.040 31.290 52.440 ;
        RECT 32.890 52.040 33.290 52.440 ;
        RECT 34.890 52.040 35.290 52.440 ;
        RECT 36.890 52.040 37.290 52.440 ;
        RECT 38.890 52.040 39.290 52.440 ;
        RECT 40.890 52.040 41.290 52.440 ;
        RECT 42.890 52.040 43.290 52.440 ;
        RECT 44.890 52.040 45.290 52.440 ;
        RECT 46.890 52.040 47.290 52.440 ;
        RECT 48.890 52.040 49.290 52.440 ;
        RECT 50.890 52.040 51.290 52.440 ;
        RECT 52.890 52.040 53.290 52.440 ;
        RECT 54.890 52.040 55.290 52.440 ;
        RECT 56.890 52.040 57.290 52.440 ;
        RECT 58.890 52.040 59.290 52.440 ;
        RECT 60.890 52.040 61.290 52.440 ;
        RECT 62.890 52.040 63.290 52.440 ;
        RECT 64.890 52.040 65.290 52.440 ;
        RECT 66.890 52.040 67.290 52.440 ;
        RECT 68.890 52.040 69.290 52.440 ;
        RECT 70.890 52.040 71.290 52.440 ;
        RECT 72.890 52.040 73.290 52.440 ;
        RECT 76.280 52.040 76.700 52.120 ;
        RECT 6.890 51.840 8.540 52.040 ;
        RECT 8.890 51.840 22.540 52.040 ;
        RECT 22.890 51.840 38.540 52.040 ;
        RECT 38.890 51.840 46.540 52.040 ;
        RECT 46.890 51.840 76.700 52.040 ;
        RECT 6.890 51.440 7.290 51.840 ;
        RECT 8.890 51.440 9.290 51.840 ;
        RECT 10.890 51.440 11.290 51.840 ;
        RECT 12.890 51.440 13.290 51.840 ;
        RECT 14.890 51.440 15.290 51.840 ;
        RECT 16.890 51.440 17.290 51.840 ;
        RECT 18.890 51.440 19.290 51.840 ;
        RECT 20.890 51.440 21.290 51.840 ;
        RECT 22.890 51.440 23.290 51.840 ;
        RECT 24.890 51.440 25.290 51.840 ;
        RECT 26.890 51.440 27.290 51.840 ;
        RECT 28.890 51.440 29.290 51.840 ;
        RECT 30.890 51.440 31.290 51.840 ;
        RECT 32.890 51.440 33.290 51.840 ;
        RECT 34.890 51.440 35.290 51.840 ;
        RECT 36.890 51.440 37.290 51.840 ;
        RECT 38.890 51.440 39.290 51.840 ;
        RECT 40.890 51.440 41.290 51.840 ;
        RECT 42.890 51.440 43.290 51.840 ;
        RECT 44.890 51.440 45.290 51.840 ;
        RECT 46.890 51.440 47.290 51.840 ;
        RECT 48.890 51.440 49.290 51.840 ;
        RECT 50.890 51.440 51.290 51.840 ;
        RECT 52.890 51.440 53.290 51.840 ;
        RECT 54.890 51.440 55.290 51.840 ;
        RECT 56.890 51.440 57.290 51.840 ;
        RECT 58.890 51.440 59.290 51.840 ;
        RECT 60.890 51.440 61.290 51.840 ;
        RECT 62.890 51.440 63.290 51.840 ;
        RECT 64.890 51.440 65.290 51.840 ;
        RECT 66.890 51.440 67.290 51.840 ;
        RECT 68.890 51.440 69.290 51.840 ;
        RECT 70.890 51.440 71.290 51.840 ;
        RECT 72.890 51.440 73.290 51.840 ;
        RECT 76.280 51.760 76.700 51.840 ;
        RECT 84.415 52.040 84.835 52.120 ;
        RECT 87.825 52.040 88.225 52.440 ;
        RECT 89.825 52.040 90.225 52.440 ;
        RECT 91.825 52.040 92.225 52.440 ;
        RECT 93.825 52.040 94.225 52.440 ;
        RECT 95.825 52.040 96.225 52.440 ;
        RECT 97.825 52.040 98.225 52.440 ;
        RECT 99.825 52.040 100.225 52.440 ;
        RECT 101.825 52.040 102.225 52.440 ;
        RECT 103.825 52.040 104.225 52.440 ;
        RECT 105.825 52.040 106.225 52.440 ;
        RECT 107.825 52.040 108.225 52.440 ;
        RECT 109.825 52.040 110.225 52.440 ;
        RECT 111.825 52.040 112.225 52.440 ;
        RECT 113.825 52.040 114.225 52.440 ;
        RECT 115.825 52.040 116.225 52.440 ;
        RECT 117.825 52.040 118.225 52.440 ;
        RECT 119.825 52.040 120.225 52.440 ;
        RECT 121.825 52.040 122.225 52.440 ;
        RECT 123.825 52.040 124.225 52.440 ;
        RECT 125.825 52.040 126.225 52.440 ;
        RECT 127.825 52.040 128.225 52.440 ;
        RECT 129.825 52.040 130.225 52.440 ;
        RECT 131.825 52.040 132.225 52.440 ;
        RECT 133.825 52.040 134.225 52.440 ;
        RECT 135.825 52.040 136.225 52.440 ;
        RECT 137.825 52.040 138.225 52.440 ;
        RECT 139.825 52.040 140.225 52.440 ;
        RECT 141.825 52.040 142.225 52.440 ;
        RECT 143.825 52.040 144.225 52.440 ;
        RECT 145.825 52.040 146.225 52.440 ;
        RECT 147.825 52.040 148.225 52.440 ;
        RECT 149.825 52.040 150.225 52.440 ;
        RECT 151.825 52.040 152.225 52.440 ;
        RECT 153.825 52.040 154.225 52.440 ;
        RECT 84.415 51.840 114.225 52.040 ;
        RECT 114.575 51.840 122.225 52.040 ;
        RECT 122.575 51.840 138.225 52.040 ;
        RECT 138.575 51.840 152.225 52.040 ;
        RECT 152.575 51.840 154.225 52.040 ;
        RECT 84.415 51.760 84.835 51.840 ;
        RECT 87.825 51.440 88.225 51.840 ;
        RECT 89.825 51.440 90.225 51.840 ;
        RECT 91.825 51.440 92.225 51.840 ;
        RECT 93.825 51.440 94.225 51.840 ;
        RECT 95.825 51.440 96.225 51.840 ;
        RECT 97.825 51.440 98.225 51.840 ;
        RECT 99.825 51.440 100.225 51.840 ;
        RECT 101.825 51.440 102.225 51.840 ;
        RECT 103.825 51.440 104.225 51.840 ;
        RECT 105.825 51.440 106.225 51.840 ;
        RECT 107.825 51.440 108.225 51.840 ;
        RECT 109.825 51.440 110.225 51.840 ;
        RECT 111.825 51.440 112.225 51.840 ;
        RECT 113.825 51.440 114.225 51.840 ;
        RECT 115.825 51.440 116.225 51.840 ;
        RECT 117.825 51.440 118.225 51.840 ;
        RECT 119.825 51.440 120.225 51.840 ;
        RECT 121.825 51.440 122.225 51.840 ;
        RECT 123.825 51.440 124.225 51.840 ;
        RECT 125.825 51.440 126.225 51.840 ;
        RECT 127.825 51.440 128.225 51.840 ;
        RECT 129.825 51.440 130.225 51.840 ;
        RECT 131.825 51.440 132.225 51.840 ;
        RECT 133.825 51.440 134.225 51.840 ;
        RECT 135.825 51.440 136.225 51.840 ;
        RECT 137.825 51.440 138.225 51.840 ;
        RECT 139.825 51.440 140.225 51.840 ;
        RECT 141.825 51.440 142.225 51.840 ;
        RECT 143.825 51.440 144.225 51.840 ;
        RECT 145.825 51.440 146.225 51.840 ;
        RECT 147.825 51.440 148.225 51.840 ;
        RECT 149.825 51.440 150.225 51.840 ;
        RECT 151.825 51.440 152.225 51.840 ;
        RECT 153.825 51.440 154.225 51.840 ;
        RECT 6.960 50.590 7.220 51.440 ;
        RECT 8.990 50.590 9.190 51.440 ;
        RECT 10.990 50.590 11.190 51.440 ;
        RECT 12.990 50.590 13.190 51.440 ;
        RECT 14.990 50.590 15.190 51.440 ;
        RECT 16.990 50.590 17.190 51.440 ;
        RECT 18.990 50.590 19.190 51.440 ;
        RECT 20.990 50.590 21.190 51.440 ;
        RECT 24.990 50.590 25.190 51.440 ;
        RECT 26.990 50.590 27.190 51.440 ;
        RECT 28.990 50.590 29.190 51.440 ;
        RECT 30.990 50.590 31.190 51.440 ;
        RECT 32.990 50.590 33.190 51.440 ;
        RECT 34.990 50.590 35.190 51.440 ;
        RECT 36.990 50.590 37.190 51.440 ;
        RECT 38.990 50.590 39.190 51.440 ;
        RECT 40.990 50.590 41.190 51.440 ;
        RECT 42.990 50.590 43.190 51.440 ;
        RECT 44.990 50.590 45.190 51.440 ;
        RECT 48.990 50.590 49.190 51.440 ;
        RECT 50.990 50.590 51.190 51.440 ;
        RECT 52.990 50.590 53.190 51.440 ;
        RECT 54.990 50.590 55.190 51.440 ;
        RECT 56.990 50.590 57.190 51.440 ;
        RECT 58.990 50.590 59.190 51.440 ;
        RECT 60.990 50.590 61.190 51.440 ;
        RECT 62.990 50.590 63.190 51.440 ;
        RECT 64.990 50.590 65.190 51.440 ;
        RECT 66.990 50.590 67.190 51.440 ;
        RECT 68.990 50.590 69.190 51.440 ;
        RECT 70.990 50.590 71.190 51.440 ;
        RECT 89.925 50.590 90.125 51.440 ;
        RECT 91.925 50.590 92.125 51.440 ;
        RECT 93.925 50.590 94.125 51.440 ;
        RECT 95.925 50.590 96.125 51.440 ;
        RECT 97.925 50.590 98.125 51.440 ;
        RECT 99.925 50.590 100.125 51.440 ;
        RECT 101.925 50.590 102.125 51.440 ;
        RECT 103.925 50.590 104.125 51.440 ;
        RECT 105.925 50.590 106.125 51.440 ;
        RECT 107.925 50.590 108.125 51.440 ;
        RECT 109.925 50.590 110.125 51.440 ;
        RECT 111.925 50.590 112.125 51.440 ;
        RECT 115.925 50.590 116.125 51.440 ;
        RECT 117.925 50.590 118.125 51.440 ;
        RECT 119.925 50.590 120.125 51.440 ;
        RECT 121.925 50.590 122.125 51.440 ;
        RECT 123.925 50.590 124.125 51.440 ;
        RECT 125.925 50.590 126.125 51.440 ;
        RECT 127.925 50.590 128.125 51.440 ;
        RECT 129.925 50.590 130.125 51.440 ;
        RECT 131.925 50.590 132.125 51.440 ;
        RECT 133.925 50.590 134.125 51.440 ;
        RECT 135.925 50.590 136.125 51.440 ;
        RECT 139.925 50.590 140.125 51.440 ;
        RECT 141.925 50.590 142.125 51.440 ;
        RECT 143.925 50.590 144.125 51.440 ;
        RECT 145.925 50.590 146.125 51.440 ;
        RECT 147.925 50.590 148.125 51.440 ;
        RECT 149.925 50.590 150.125 51.440 ;
        RECT 151.925 50.590 152.125 51.440 ;
        RECT 153.895 50.590 154.155 51.440 ;
        RECT 6.890 50.190 7.290 50.590 ;
        RECT 8.890 50.190 9.290 50.590 ;
        RECT 10.890 50.190 11.290 50.590 ;
        RECT 12.890 50.190 13.290 50.590 ;
        RECT 14.890 50.190 15.290 50.590 ;
        RECT 16.890 50.190 17.290 50.590 ;
        RECT 18.890 50.190 19.290 50.590 ;
        RECT 20.890 50.190 21.290 50.590 ;
        RECT 22.890 50.190 23.290 50.590 ;
        RECT 24.890 50.190 25.290 50.590 ;
        RECT 26.890 50.190 27.290 50.590 ;
        RECT 28.890 50.190 29.290 50.590 ;
        RECT 30.890 50.190 31.290 50.590 ;
        RECT 32.890 50.190 33.290 50.590 ;
        RECT 34.890 50.190 35.290 50.590 ;
        RECT 36.890 50.190 37.290 50.590 ;
        RECT 38.890 50.190 39.290 50.590 ;
        RECT 40.890 50.190 41.290 50.590 ;
        RECT 42.890 50.190 43.290 50.590 ;
        RECT 44.890 50.190 45.290 50.590 ;
        RECT 46.890 50.190 47.290 50.590 ;
        RECT 48.890 50.190 49.290 50.590 ;
        RECT 50.890 50.190 51.290 50.590 ;
        RECT 52.890 50.190 53.290 50.590 ;
        RECT 54.890 50.190 55.290 50.590 ;
        RECT 56.890 50.190 57.290 50.590 ;
        RECT 58.890 50.190 59.290 50.590 ;
        RECT 60.890 50.190 61.290 50.590 ;
        RECT 62.890 50.190 63.290 50.590 ;
        RECT 64.890 50.190 65.290 50.590 ;
        RECT 66.890 50.190 67.290 50.590 ;
        RECT 68.890 50.190 69.290 50.590 ;
        RECT 70.890 50.190 71.290 50.590 ;
        RECT 72.890 50.190 73.290 50.590 ;
        RECT 87.825 50.190 88.225 50.590 ;
        RECT 89.825 50.190 90.225 50.590 ;
        RECT 91.825 50.190 92.225 50.590 ;
        RECT 93.825 50.190 94.225 50.590 ;
        RECT 95.825 50.190 96.225 50.590 ;
        RECT 97.825 50.190 98.225 50.590 ;
        RECT 99.825 50.190 100.225 50.590 ;
        RECT 101.825 50.190 102.225 50.590 ;
        RECT 103.825 50.190 104.225 50.590 ;
        RECT 105.825 50.190 106.225 50.590 ;
        RECT 107.825 50.190 108.225 50.590 ;
        RECT 109.825 50.190 110.225 50.590 ;
        RECT 111.825 50.190 112.225 50.590 ;
        RECT 113.825 50.190 114.225 50.590 ;
        RECT 115.825 50.190 116.225 50.590 ;
        RECT 117.825 50.190 118.225 50.590 ;
        RECT 119.825 50.190 120.225 50.590 ;
        RECT 121.825 50.190 122.225 50.590 ;
        RECT 123.825 50.190 124.225 50.590 ;
        RECT 125.825 50.190 126.225 50.590 ;
        RECT 127.825 50.190 128.225 50.590 ;
        RECT 129.825 50.190 130.225 50.590 ;
        RECT 131.825 50.190 132.225 50.590 ;
        RECT 133.825 50.190 134.225 50.590 ;
        RECT 135.825 50.190 136.225 50.590 ;
        RECT 137.825 50.190 138.225 50.590 ;
        RECT 139.825 50.190 140.225 50.590 ;
        RECT 141.825 50.190 142.225 50.590 ;
        RECT 143.825 50.190 144.225 50.590 ;
        RECT 145.825 50.190 146.225 50.590 ;
        RECT 147.825 50.190 148.225 50.590 ;
        RECT 149.825 50.190 150.225 50.590 ;
        RECT 151.825 50.190 152.225 50.590 ;
        RECT 153.825 50.190 154.225 50.590 ;
        RECT 6.890 49.990 8.540 50.190 ;
        RECT 8.890 49.990 24.540 50.190 ;
        RECT 24.890 49.990 38.540 50.190 ;
        RECT 38.890 49.990 48.540 50.190 ;
        RECT 48.890 49.990 74.540 50.190 ;
        RECT 86.575 49.990 112.225 50.190 ;
        RECT 112.575 49.990 122.225 50.190 ;
        RECT 122.575 49.990 136.225 50.190 ;
        RECT 136.575 49.990 152.225 50.190 ;
        RECT 152.575 49.990 154.225 50.190 ;
        RECT 6.890 49.590 7.290 49.990 ;
        RECT 8.890 49.590 9.290 49.990 ;
        RECT 10.890 49.590 11.290 49.990 ;
        RECT 12.890 49.590 13.290 49.990 ;
        RECT 14.890 49.590 15.290 49.990 ;
        RECT 16.890 49.590 17.290 49.990 ;
        RECT 18.890 49.590 19.290 49.990 ;
        RECT 20.890 49.590 21.290 49.990 ;
        RECT 22.890 49.590 23.290 49.990 ;
        RECT 24.890 49.590 25.290 49.990 ;
        RECT 26.890 49.590 27.290 49.990 ;
        RECT 28.890 49.590 29.290 49.990 ;
        RECT 30.890 49.590 31.290 49.990 ;
        RECT 32.890 49.590 33.290 49.990 ;
        RECT 34.890 49.590 35.290 49.990 ;
        RECT 36.890 49.590 37.290 49.990 ;
        RECT 38.890 49.590 39.290 49.990 ;
        RECT 40.890 49.590 41.290 49.990 ;
        RECT 42.890 49.590 43.290 49.990 ;
        RECT 44.890 49.590 45.290 49.990 ;
        RECT 46.890 49.590 47.290 49.990 ;
        RECT 48.890 49.590 49.290 49.990 ;
        RECT 50.890 49.590 51.290 49.990 ;
        RECT 52.890 49.590 53.290 49.990 ;
        RECT 54.890 49.590 55.290 49.990 ;
        RECT 56.890 49.590 57.290 49.990 ;
        RECT 58.890 49.590 59.290 49.990 ;
        RECT 60.890 49.590 61.290 49.990 ;
        RECT 62.890 49.590 63.290 49.990 ;
        RECT 64.890 49.590 65.290 49.990 ;
        RECT 66.890 49.590 67.290 49.990 ;
        RECT 68.890 49.590 69.290 49.990 ;
        RECT 70.890 49.590 71.290 49.990 ;
        RECT 72.890 49.590 73.290 49.990 ;
        RECT 87.825 49.590 88.225 49.990 ;
        RECT 89.825 49.590 90.225 49.990 ;
        RECT 91.825 49.590 92.225 49.990 ;
        RECT 93.825 49.590 94.225 49.990 ;
        RECT 95.825 49.590 96.225 49.990 ;
        RECT 97.825 49.590 98.225 49.990 ;
        RECT 99.825 49.590 100.225 49.990 ;
        RECT 101.825 49.590 102.225 49.990 ;
        RECT 103.825 49.590 104.225 49.990 ;
        RECT 105.825 49.590 106.225 49.990 ;
        RECT 107.825 49.590 108.225 49.990 ;
        RECT 109.825 49.590 110.225 49.990 ;
        RECT 111.825 49.590 112.225 49.990 ;
        RECT 113.825 49.590 114.225 49.990 ;
        RECT 115.825 49.590 116.225 49.990 ;
        RECT 117.825 49.590 118.225 49.990 ;
        RECT 119.825 49.590 120.225 49.990 ;
        RECT 121.825 49.590 122.225 49.990 ;
        RECT 123.825 49.590 124.225 49.990 ;
        RECT 125.825 49.590 126.225 49.990 ;
        RECT 127.825 49.590 128.225 49.990 ;
        RECT 129.825 49.590 130.225 49.990 ;
        RECT 131.825 49.590 132.225 49.990 ;
        RECT 133.825 49.590 134.225 49.990 ;
        RECT 135.825 49.590 136.225 49.990 ;
        RECT 137.825 49.590 138.225 49.990 ;
        RECT 139.825 49.590 140.225 49.990 ;
        RECT 141.825 49.590 142.225 49.990 ;
        RECT 143.825 49.590 144.225 49.990 ;
        RECT 145.825 49.590 146.225 49.990 ;
        RECT 147.825 49.590 148.225 49.990 ;
        RECT 149.825 49.590 150.225 49.990 ;
        RECT 151.825 49.590 152.225 49.990 ;
        RECT 153.825 49.590 154.225 49.990 ;
        RECT 6.960 48.740 7.220 49.590 ;
        RECT 8.990 48.740 9.190 49.590 ;
        RECT 10.990 48.740 11.190 49.590 ;
        RECT 12.990 48.740 13.190 49.590 ;
        RECT 14.990 48.740 15.190 49.590 ;
        RECT 16.990 48.740 17.190 49.590 ;
        RECT 18.990 48.740 19.190 49.590 ;
        RECT 20.990 48.740 21.190 49.590 ;
        RECT 22.990 48.740 23.190 49.590 ;
        RECT 24.990 48.740 25.190 49.590 ;
        RECT 26.990 48.740 27.190 49.590 ;
        RECT 28.990 48.740 29.190 49.590 ;
        RECT 30.990 48.740 31.190 49.590 ;
        RECT 32.990 48.740 33.190 49.590 ;
        RECT 34.990 48.740 35.190 49.590 ;
        RECT 36.990 48.740 37.190 49.590 ;
        RECT 38.990 48.740 39.190 49.590 ;
        RECT 40.990 48.740 41.190 49.590 ;
        RECT 42.990 48.740 43.190 49.590 ;
        RECT 44.990 48.740 45.190 49.590 ;
        RECT 46.990 48.740 47.190 49.590 ;
        RECT 48.990 48.740 49.190 49.590 ;
        RECT 50.990 48.740 51.190 49.590 ;
        RECT 52.990 48.740 53.190 49.590 ;
        RECT 54.990 48.740 55.190 49.590 ;
        RECT 56.990 48.740 57.190 49.590 ;
        RECT 58.990 48.740 59.190 49.590 ;
        RECT 60.990 48.740 61.190 49.590 ;
        RECT 62.990 48.740 63.190 49.590 ;
        RECT 64.990 48.740 65.190 49.590 ;
        RECT 66.990 48.740 67.190 49.590 ;
        RECT 68.990 48.740 69.190 49.590 ;
        RECT 70.990 48.740 71.190 49.590 ;
        RECT 89.925 48.740 90.125 49.590 ;
        RECT 91.925 48.740 92.125 49.590 ;
        RECT 93.925 48.740 94.125 49.590 ;
        RECT 95.925 48.740 96.125 49.590 ;
        RECT 97.925 48.740 98.125 49.590 ;
        RECT 99.925 48.740 100.125 49.590 ;
        RECT 101.925 48.740 102.125 49.590 ;
        RECT 103.925 48.740 104.125 49.590 ;
        RECT 105.925 48.740 106.125 49.590 ;
        RECT 107.925 48.740 108.125 49.590 ;
        RECT 109.925 48.740 110.125 49.590 ;
        RECT 111.925 48.740 112.125 49.590 ;
        RECT 113.925 48.740 114.125 49.590 ;
        RECT 115.925 48.740 116.125 49.590 ;
        RECT 117.925 48.740 118.125 49.590 ;
        RECT 119.925 48.740 120.125 49.590 ;
        RECT 121.925 48.740 122.125 49.590 ;
        RECT 123.925 48.740 124.125 49.590 ;
        RECT 125.925 48.740 126.125 49.590 ;
        RECT 127.925 48.740 128.125 49.590 ;
        RECT 129.925 48.740 130.125 49.590 ;
        RECT 131.925 48.740 132.125 49.590 ;
        RECT 133.925 48.740 134.125 49.590 ;
        RECT 135.925 48.740 136.125 49.590 ;
        RECT 137.925 48.740 138.125 49.590 ;
        RECT 139.925 48.740 140.125 49.590 ;
        RECT 141.925 48.740 142.125 49.590 ;
        RECT 143.925 48.740 144.125 49.590 ;
        RECT 145.925 48.740 146.125 49.590 ;
        RECT 147.925 48.740 148.125 49.590 ;
        RECT 149.925 48.740 150.125 49.590 ;
        RECT 151.925 48.740 152.125 49.590 ;
        RECT 153.895 48.740 154.155 49.590 ;
        RECT 6.890 48.340 7.290 48.740 ;
        RECT 8.890 48.340 9.290 48.740 ;
        RECT 10.890 48.340 11.290 48.740 ;
        RECT 12.890 48.340 13.290 48.740 ;
        RECT 14.890 48.340 15.290 48.740 ;
        RECT 16.890 48.340 17.290 48.740 ;
        RECT 18.890 48.340 19.290 48.740 ;
        RECT 20.890 48.340 21.290 48.740 ;
        RECT 22.890 48.340 23.290 48.740 ;
        RECT 24.890 48.340 25.290 48.740 ;
        RECT 26.890 48.340 27.290 48.740 ;
        RECT 28.890 48.340 29.290 48.740 ;
        RECT 30.890 48.340 31.290 48.740 ;
        RECT 32.890 48.340 33.290 48.740 ;
        RECT 34.890 48.340 35.290 48.740 ;
        RECT 36.890 48.340 37.290 48.740 ;
        RECT 38.890 48.340 39.290 48.740 ;
        RECT 40.890 48.340 41.290 48.740 ;
        RECT 42.890 48.340 43.290 48.740 ;
        RECT 44.890 48.340 45.290 48.740 ;
        RECT 46.890 48.340 47.290 48.740 ;
        RECT 48.890 48.340 49.290 48.740 ;
        RECT 50.890 48.340 51.290 48.740 ;
        RECT 52.890 48.340 53.290 48.740 ;
        RECT 54.890 48.340 55.290 48.740 ;
        RECT 56.890 48.340 57.290 48.740 ;
        RECT 58.890 48.340 59.290 48.740 ;
        RECT 60.890 48.340 61.290 48.740 ;
        RECT 62.890 48.340 63.290 48.740 ;
        RECT 64.890 48.340 65.290 48.740 ;
        RECT 66.890 48.340 67.290 48.740 ;
        RECT 68.890 48.340 69.290 48.740 ;
        RECT 70.890 48.340 71.290 48.740 ;
        RECT 72.890 48.340 73.290 48.740 ;
        RECT 87.825 48.340 88.225 48.740 ;
        RECT 89.825 48.340 90.225 48.740 ;
        RECT 91.825 48.340 92.225 48.740 ;
        RECT 93.825 48.340 94.225 48.740 ;
        RECT 95.825 48.340 96.225 48.740 ;
        RECT 97.825 48.340 98.225 48.740 ;
        RECT 99.825 48.340 100.225 48.740 ;
        RECT 101.825 48.340 102.225 48.740 ;
        RECT 103.825 48.340 104.225 48.740 ;
        RECT 105.825 48.340 106.225 48.740 ;
        RECT 107.825 48.340 108.225 48.740 ;
        RECT 109.825 48.340 110.225 48.740 ;
        RECT 111.825 48.340 112.225 48.740 ;
        RECT 113.825 48.340 114.225 48.740 ;
        RECT 115.825 48.340 116.225 48.740 ;
        RECT 117.825 48.340 118.225 48.740 ;
        RECT 119.825 48.340 120.225 48.740 ;
        RECT 121.825 48.340 122.225 48.740 ;
        RECT 123.825 48.340 124.225 48.740 ;
        RECT 125.825 48.340 126.225 48.740 ;
        RECT 127.825 48.340 128.225 48.740 ;
        RECT 129.825 48.340 130.225 48.740 ;
        RECT 131.825 48.340 132.225 48.740 ;
        RECT 133.825 48.340 134.225 48.740 ;
        RECT 135.825 48.340 136.225 48.740 ;
        RECT 137.825 48.340 138.225 48.740 ;
        RECT 139.825 48.340 140.225 48.740 ;
        RECT 141.825 48.340 142.225 48.740 ;
        RECT 143.825 48.340 144.225 48.740 ;
        RECT 145.825 48.340 146.225 48.740 ;
        RECT 147.825 48.340 148.225 48.740 ;
        RECT 149.825 48.340 150.225 48.740 ;
        RECT 151.825 48.340 152.225 48.740 ;
        RECT 153.825 48.340 154.225 48.740 ;
        RECT 6.890 48.140 8.540 48.340 ;
        RECT 8.890 48.140 24.540 48.340 ;
        RECT 24.890 48.140 38.540 48.340 ;
        RECT 38.890 48.140 48.540 48.340 ;
        RECT 48.890 48.140 74.540 48.340 ;
        RECT 86.575 48.140 112.225 48.340 ;
        RECT 112.575 48.140 122.225 48.340 ;
        RECT 122.575 48.140 136.225 48.340 ;
        RECT 136.575 48.140 152.225 48.340 ;
        RECT 152.575 48.140 154.225 48.340 ;
        RECT 6.890 47.740 7.290 48.140 ;
        RECT 8.890 47.740 9.290 48.140 ;
        RECT 10.890 47.740 11.290 48.140 ;
        RECT 12.890 47.740 13.290 48.140 ;
        RECT 14.890 47.740 15.290 48.140 ;
        RECT 16.890 47.740 17.290 48.140 ;
        RECT 18.890 47.740 19.290 48.140 ;
        RECT 20.890 47.740 21.290 48.140 ;
        RECT 22.890 47.740 23.290 48.140 ;
        RECT 24.890 47.740 25.290 48.140 ;
        RECT 26.890 47.740 27.290 48.140 ;
        RECT 28.890 47.740 29.290 48.140 ;
        RECT 30.890 47.740 31.290 48.140 ;
        RECT 32.890 47.740 33.290 48.140 ;
        RECT 34.890 47.740 35.290 48.140 ;
        RECT 36.890 47.740 37.290 48.140 ;
        RECT 38.890 47.740 39.290 48.140 ;
        RECT 40.890 47.740 41.290 48.140 ;
        RECT 42.890 47.740 43.290 48.140 ;
        RECT 44.890 47.740 45.290 48.140 ;
        RECT 46.890 47.740 47.290 48.140 ;
        RECT 48.890 47.740 49.290 48.140 ;
        RECT 50.890 47.740 51.290 48.140 ;
        RECT 52.890 47.740 53.290 48.140 ;
        RECT 54.890 47.740 55.290 48.140 ;
        RECT 56.890 47.740 57.290 48.140 ;
        RECT 58.890 47.740 59.290 48.140 ;
        RECT 60.890 47.740 61.290 48.140 ;
        RECT 62.890 47.740 63.290 48.140 ;
        RECT 64.890 47.740 65.290 48.140 ;
        RECT 66.890 47.740 67.290 48.140 ;
        RECT 68.890 47.740 69.290 48.140 ;
        RECT 70.890 47.740 71.290 48.140 ;
        RECT 72.890 47.740 73.290 48.140 ;
        RECT 87.825 47.740 88.225 48.140 ;
        RECT 89.825 47.740 90.225 48.140 ;
        RECT 91.825 47.740 92.225 48.140 ;
        RECT 93.825 47.740 94.225 48.140 ;
        RECT 95.825 47.740 96.225 48.140 ;
        RECT 97.825 47.740 98.225 48.140 ;
        RECT 99.825 47.740 100.225 48.140 ;
        RECT 101.825 47.740 102.225 48.140 ;
        RECT 103.825 47.740 104.225 48.140 ;
        RECT 105.825 47.740 106.225 48.140 ;
        RECT 107.825 47.740 108.225 48.140 ;
        RECT 109.825 47.740 110.225 48.140 ;
        RECT 111.825 47.740 112.225 48.140 ;
        RECT 113.825 47.740 114.225 48.140 ;
        RECT 115.825 47.740 116.225 48.140 ;
        RECT 117.825 47.740 118.225 48.140 ;
        RECT 119.825 47.740 120.225 48.140 ;
        RECT 121.825 47.740 122.225 48.140 ;
        RECT 123.825 47.740 124.225 48.140 ;
        RECT 125.825 47.740 126.225 48.140 ;
        RECT 127.825 47.740 128.225 48.140 ;
        RECT 129.825 47.740 130.225 48.140 ;
        RECT 131.825 47.740 132.225 48.140 ;
        RECT 133.825 47.740 134.225 48.140 ;
        RECT 135.825 47.740 136.225 48.140 ;
        RECT 137.825 47.740 138.225 48.140 ;
        RECT 139.825 47.740 140.225 48.140 ;
        RECT 141.825 47.740 142.225 48.140 ;
        RECT 143.825 47.740 144.225 48.140 ;
        RECT 145.825 47.740 146.225 48.140 ;
        RECT 147.825 47.740 148.225 48.140 ;
        RECT 149.825 47.740 150.225 48.140 ;
        RECT 151.825 47.740 152.225 48.140 ;
        RECT 153.825 47.740 154.225 48.140 ;
        RECT 6.960 46.890 7.220 47.740 ;
        RECT 8.990 46.890 9.190 47.740 ;
        RECT 10.990 46.890 11.190 47.740 ;
        RECT 12.990 46.890 13.190 47.740 ;
        RECT 14.990 46.890 15.190 47.740 ;
        RECT 16.990 46.890 17.190 47.740 ;
        RECT 18.990 46.890 19.190 47.740 ;
        RECT 20.990 46.890 21.190 47.740 ;
        RECT 22.990 46.890 23.190 47.740 ;
        RECT 24.990 46.890 25.190 47.740 ;
        RECT 26.990 46.890 27.190 47.740 ;
        RECT 28.990 46.890 29.190 47.740 ;
        RECT 30.990 46.890 31.190 47.740 ;
        RECT 32.990 46.890 33.190 47.740 ;
        RECT 34.990 46.890 35.190 47.740 ;
        RECT 36.990 46.890 37.190 47.740 ;
        RECT 38.990 46.890 39.190 47.740 ;
        RECT 40.990 46.890 41.190 47.740 ;
        RECT 42.990 46.890 43.190 47.740 ;
        RECT 44.990 46.890 45.190 47.740 ;
        RECT 46.990 46.890 47.190 47.740 ;
        RECT 113.925 46.890 114.125 47.740 ;
        RECT 115.925 46.890 116.125 47.740 ;
        RECT 117.925 46.890 118.125 47.740 ;
        RECT 119.925 46.890 120.125 47.740 ;
        RECT 121.925 46.890 122.125 47.740 ;
        RECT 123.925 46.890 124.125 47.740 ;
        RECT 125.925 46.890 126.125 47.740 ;
        RECT 127.925 46.890 128.125 47.740 ;
        RECT 129.925 46.890 130.125 47.740 ;
        RECT 131.925 46.890 132.125 47.740 ;
        RECT 133.925 46.890 134.125 47.740 ;
        RECT 135.925 46.890 136.125 47.740 ;
        RECT 137.925 46.890 138.125 47.740 ;
        RECT 139.925 46.890 140.125 47.740 ;
        RECT 141.925 46.890 142.125 47.740 ;
        RECT 143.925 46.890 144.125 47.740 ;
        RECT 145.925 46.890 146.125 47.740 ;
        RECT 147.925 46.890 148.125 47.740 ;
        RECT 149.925 46.890 150.125 47.740 ;
        RECT 151.925 46.890 152.125 47.740 ;
        RECT 153.895 46.890 154.155 47.740 ;
        RECT 6.890 46.490 7.290 46.890 ;
        RECT 8.890 46.490 9.290 46.890 ;
        RECT 10.890 46.490 11.290 46.890 ;
        RECT 12.890 46.490 13.290 46.890 ;
        RECT 14.890 46.490 15.290 46.890 ;
        RECT 16.890 46.490 17.290 46.890 ;
        RECT 18.890 46.490 19.290 46.890 ;
        RECT 20.890 46.490 21.290 46.890 ;
        RECT 22.890 46.490 23.290 46.890 ;
        RECT 24.890 46.490 25.290 46.890 ;
        RECT 26.890 46.490 27.290 46.890 ;
        RECT 28.890 46.490 29.290 46.890 ;
        RECT 30.890 46.490 31.290 46.890 ;
        RECT 32.890 46.490 33.290 46.890 ;
        RECT 34.890 46.490 35.290 46.890 ;
        RECT 36.890 46.490 37.290 46.890 ;
        RECT 38.890 46.490 39.290 46.890 ;
        RECT 40.890 46.490 41.290 46.890 ;
        RECT 42.890 46.490 43.290 46.890 ;
        RECT 44.890 46.490 45.290 46.890 ;
        RECT 46.890 46.490 47.290 46.890 ;
        RECT 48.890 46.490 49.290 46.890 ;
        RECT 50.890 46.490 51.290 46.890 ;
        RECT 52.890 46.490 53.290 46.890 ;
        RECT 54.890 46.490 55.290 46.890 ;
        RECT 56.890 46.490 57.290 46.890 ;
        RECT 58.890 46.490 59.290 46.890 ;
        RECT 60.890 46.490 61.290 46.890 ;
        RECT 62.890 46.490 63.290 46.890 ;
        RECT 64.890 46.490 65.290 46.890 ;
        RECT 66.890 46.490 67.290 46.890 ;
        RECT 68.890 46.490 69.290 46.890 ;
        RECT 70.890 46.490 71.290 46.890 ;
        RECT 72.890 46.490 73.290 46.890 ;
        RECT 75.830 46.490 76.250 46.570 ;
        RECT 6.890 46.290 8.540 46.490 ;
        RECT 8.890 46.290 24.540 46.490 ;
        RECT 24.890 46.290 38.540 46.490 ;
        RECT 38.890 46.290 76.250 46.490 ;
        RECT 6.890 45.890 7.290 46.290 ;
        RECT 8.890 45.890 9.290 46.290 ;
        RECT 10.890 45.890 11.290 46.290 ;
        RECT 12.890 45.890 13.290 46.290 ;
        RECT 14.890 45.890 15.290 46.290 ;
        RECT 16.890 45.890 17.290 46.290 ;
        RECT 18.890 45.890 19.290 46.290 ;
        RECT 20.890 45.890 21.290 46.290 ;
        RECT 22.890 45.890 23.290 46.290 ;
        RECT 24.890 45.890 25.290 46.290 ;
        RECT 26.890 45.890 27.290 46.290 ;
        RECT 28.890 45.890 29.290 46.290 ;
        RECT 30.890 45.890 31.290 46.290 ;
        RECT 32.890 45.890 33.290 46.290 ;
        RECT 34.890 45.890 35.290 46.290 ;
        RECT 36.890 45.890 37.290 46.290 ;
        RECT 38.890 45.890 39.290 46.290 ;
        RECT 40.890 45.890 41.290 46.290 ;
        RECT 42.890 45.890 43.290 46.290 ;
        RECT 44.890 45.890 45.290 46.290 ;
        RECT 46.890 45.890 47.290 46.290 ;
        RECT 48.890 45.890 49.290 46.290 ;
        RECT 50.890 45.890 51.290 46.290 ;
        RECT 52.890 45.890 53.290 46.290 ;
        RECT 54.890 45.890 55.290 46.290 ;
        RECT 56.890 45.890 57.290 46.290 ;
        RECT 58.890 45.890 59.290 46.290 ;
        RECT 60.890 45.890 61.290 46.290 ;
        RECT 62.890 45.890 63.290 46.290 ;
        RECT 64.890 45.890 65.290 46.290 ;
        RECT 66.890 45.890 67.290 46.290 ;
        RECT 68.890 45.890 69.290 46.290 ;
        RECT 70.890 45.890 71.290 46.290 ;
        RECT 72.890 45.890 73.290 46.290 ;
        RECT 75.830 46.210 76.250 46.290 ;
        RECT 84.865 46.490 85.285 46.570 ;
        RECT 87.825 46.490 88.225 46.890 ;
        RECT 89.825 46.490 90.225 46.890 ;
        RECT 91.825 46.490 92.225 46.890 ;
        RECT 93.825 46.490 94.225 46.890 ;
        RECT 95.825 46.490 96.225 46.890 ;
        RECT 97.825 46.490 98.225 46.890 ;
        RECT 99.825 46.490 100.225 46.890 ;
        RECT 101.825 46.490 102.225 46.890 ;
        RECT 103.825 46.490 104.225 46.890 ;
        RECT 105.825 46.490 106.225 46.890 ;
        RECT 107.825 46.490 108.225 46.890 ;
        RECT 109.825 46.490 110.225 46.890 ;
        RECT 111.825 46.490 112.225 46.890 ;
        RECT 113.825 46.490 114.225 46.890 ;
        RECT 115.825 46.490 116.225 46.890 ;
        RECT 117.825 46.490 118.225 46.890 ;
        RECT 119.825 46.490 120.225 46.890 ;
        RECT 121.825 46.490 122.225 46.890 ;
        RECT 123.825 46.490 124.225 46.890 ;
        RECT 125.825 46.490 126.225 46.890 ;
        RECT 127.825 46.490 128.225 46.890 ;
        RECT 129.825 46.490 130.225 46.890 ;
        RECT 131.825 46.490 132.225 46.890 ;
        RECT 133.825 46.490 134.225 46.890 ;
        RECT 135.825 46.490 136.225 46.890 ;
        RECT 137.825 46.490 138.225 46.890 ;
        RECT 139.825 46.490 140.225 46.890 ;
        RECT 141.825 46.490 142.225 46.890 ;
        RECT 143.825 46.490 144.225 46.890 ;
        RECT 145.825 46.490 146.225 46.890 ;
        RECT 147.825 46.490 148.225 46.890 ;
        RECT 149.825 46.490 150.225 46.890 ;
        RECT 151.825 46.490 152.225 46.890 ;
        RECT 153.825 46.490 154.225 46.890 ;
        RECT 84.865 46.290 122.225 46.490 ;
        RECT 122.575 46.290 136.225 46.490 ;
        RECT 136.575 46.290 152.225 46.490 ;
        RECT 152.575 46.290 154.225 46.490 ;
        RECT 84.865 46.210 85.285 46.290 ;
        RECT 87.825 45.890 88.225 46.290 ;
        RECT 89.825 45.890 90.225 46.290 ;
        RECT 91.825 45.890 92.225 46.290 ;
        RECT 93.825 45.890 94.225 46.290 ;
        RECT 95.825 45.890 96.225 46.290 ;
        RECT 97.825 45.890 98.225 46.290 ;
        RECT 99.825 45.890 100.225 46.290 ;
        RECT 101.825 45.890 102.225 46.290 ;
        RECT 103.825 45.890 104.225 46.290 ;
        RECT 105.825 45.890 106.225 46.290 ;
        RECT 107.825 45.890 108.225 46.290 ;
        RECT 109.825 45.890 110.225 46.290 ;
        RECT 111.825 45.890 112.225 46.290 ;
        RECT 113.825 45.890 114.225 46.290 ;
        RECT 115.825 45.890 116.225 46.290 ;
        RECT 117.825 45.890 118.225 46.290 ;
        RECT 119.825 45.890 120.225 46.290 ;
        RECT 121.825 45.890 122.225 46.290 ;
        RECT 123.825 45.890 124.225 46.290 ;
        RECT 125.825 45.890 126.225 46.290 ;
        RECT 127.825 45.890 128.225 46.290 ;
        RECT 129.825 45.890 130.225 46.290 ;
        RECT 131.825 45.890 132.225 46.290 ;
        RECT 133.825 45.890 134.225 46.290 ;
        RECT 135.825 45.890 136.225 46.290 ;
        RECT 137.825 45.890 138.225 46.290 ;
        RECT 139.825 45.890 140.225 46.290 ;
        RECT 141.825 45.890 142.225 46.290 ;
        RECT 143.825 45.890 144.225 46.290 ;
        RECT 145.825 45.890 146.225 46.290 ;
        RECT 147.825 45.890 148.225 46.290 ;
        RECT 149.825 45.890 150.225 46.290 ;
        RECT 151.825 45.890 152.225 46.290 ;
        RECT 153.825 45.890 154.225 46.290 ;
        RECT 6.960 45.040 7.220 45.890 ;
        RECT 8.990 45.040 9.190 45.890 ;
        RECT 10.990 45.040 11.190 45.890 ;
        RECT 12.990 45.040 13.190 45.890 ;
        RECT 14.990 45.040 15.190 45.890 ;
        RECT 16.990 45.040 17.190 45.890 ;
        RECT 18.990 45.040 19.190 45.890 ;
        RECT 20.990 45.040 21.190 45.890 ;
        RECT 22.990 45.040 23.190 45.890 ;
        RECT 24.990 45.040 25.190 45.890 ;
        RECT 26.990 45.040 27.190 45.890 ;
        RECT 28.990 45.040 29.190 45.890 ;
        RECT 30.990 45.040 31.190 45.890 ;
        RECT 32.990 45.040 33.190 45.890 ;
        RECT 34.990 45.040 35.190 45.890 ;
        RECT 36.990 45.040 37.190 45.890 ;
        RECT 38.990 45.040 39.190 45.890 ;
        RECT 40.990 45.040 41.190 45.890 ;
        RECT 42.990 45.040 43.190 45.890 ;
        RECT 44.990 45.040 45.190 45.890 ;
        RECT 46.990 45.040 47.190 45.890 ;
        RECT 48.990 45.040 49.190 45.890 ;
        RECT 50.990 45.040 51.190 45.890 ;
        RECT 52.990 45.040 53.190 45.890 ;
        RECT 54.990 45.040 55.190 45.890 ;
        RECT 56.990 45.040 57.190 45.890 ;
        RECT 58.990 45.040 59.190 45.890 ;
        RECT 60.990 45.040 61.190 45.890 ;
        RECT 62.990 45.040 63.190 45.890 ;
        RECT 64.990 45.040 65.190 45.890 ;
        RECT 66.990 45.040 67.190 45.890 ;
        RECT 68.990 45.040 69.190 45.890 ;
        RECT 70.990 45.040 71.190 45.890 ;
        RECT 89.925 45.040 90.125 45.890 ;
        RECT 91.925 45.040 92.125 45.890 ;
        RECT 93.925 45.040 94.125 45.890 ;
        RECT 95.925 45.040 96.125 45.890 ;
        RECT 97.925 45.040 98.125 45.890 ;
        RECT 99.925 45.040 100.125 45.890 ;
        RECT 101.925 45.040 102.125 45.890 ;
        RECT 103.925 45.040 104.125 45.890 ;
        RECT 105.925 45.040 106.125 45.890 ;
        RECT 107.925 45.040 108.125 45.890 ;
        RECT 109.925 45.040 110.125 45.890 ;
        RECT 111.925 45.040 112.125 45.890 ;
        RECT 113.925 45.040 114.125 45.890 ;
        RECT 115.925 45.040 116.125 45.890 ;
        RECT 117.925 45.040 118.125 45.890 ;
        RECT 119.925 45.040 120.125 45.890 ;
        RECT 121.925 45.040 122.125 45.890 ;
        RECT 123.925 45.040 124.125 45.890 ;
        RECT 125.925 45.040 126.125 45.890 ;
        RECT 127.925 45.040 128.125 45.890 ;
        RECT 129.925 45.040 130.125 45.890 ;
        RECT 131.925 45.040 132.125 45.890 ;
        RECT 133.925 45.040 134.125 45.890 ;
        RECT 135.925 45.040 136.125 45.890 ;
        RECT 137.925 45.040 138.125 45.890 ;
        RECT 139.925 45.040 140.125 45.890 ;
        RECT 141.925 45.040 142.125 45.890 ;
        RECT 143.925 45.040 144.125 45.890 ;
        RECT 145.925 45.040 146.125 45.890 ;
        RECT 147.925 45.040 148.125 45.890 ;
        RECT 149.925 45.040 150.125 45.890 ;
        RECT 151.925 45.040 152.125 45.890 ;
        RECT 153.895 45.040 154.155 45.890 ;
        RECT 6.890 44.640 7.290 45.040 ;
        RECT 8.890 44.640 9.290 45.040 ;
        RECT 10.890 44.640 11.290 45.040 ;
        RECT 12.890 44.640 13.290 45.040 ;
        RECT 14.890 44.640 15.290 45.040 ;
        RECT 16.890 44.640 17.290 45.040 ;
        RECT 18.890 44.640 19.290 45.040 ;
        RECT 20.890 44.640 21.290 45.040 ;
        RECT 22.890 44.640 23.290 45.040 ;
        RECT 24.890 44.640 25.290 45.040 ;
        RECT 26.890 44.640 27.290 45.040 ;
        RECT 28.890 44.640 29.290 45.040 ;
        RECT 30.890 44.640 31.290 45.040 ;
        RECT 32.890 44.640 33.290 45.040 ;
        RECT 34.890 44.640 35.290 45.040 ;
        RECT 36.890 44.640 37.290 45.040 ;
        RECT 38.890 44.640 39.290 45.040 ;
        RECT 40.890 44.640 41.290 45.040 ;
        RECT 42.890 44.640 43.290 45.040 ;
        RECT 44.890 44.640 45.290 45.040 ;
        RECT 46.890 44.640 47.290 45.040 ;
        RECT 48.890 44.640 49.290 45.040 ;
        RECT 50.890 44.640 51.290 45.040 ;
        RECT 52.890 44.640 53.290 45.040 ;
        RECT 54.890 44.640 55.290 45.040 ;
        RECT 56.890 44.640 57.290 45.040 ;
        RECT 58.890 44.640 59.290 45.040 ;
        RECT 60.890 44.640 61.290 45.040 ;
        RECT 62.890 44.640 63.290 45.040 ;
        RECT 64.890 44.640 65.290 45.040 ;
        RECT 66.890 44.640 67.290 45.040 ;
        RECT 68.890 44.640 69.290 45.040 ;
        RECT 70.890 44.640 71.290 45.040 ;
        RECT 72.890 44.640 73.290 45.040 ;
        RECT 87.825 44.640 88.225 45.040 ;
        RECT 89.825 44.640 90.225 45.040 ;
        RECT 91.825 44.640 92.225 45.040 ;
        RECT 93.825 44.640 94.225 45.040 ;
        RECT 95.825 44.640 96.225 45.040 ;
        RECT 97.825 44.640 98.225 45.040 ;
        RECT 99.825 44.640 100.225 45.040 ;
        RECT 101.825 44.640 102.225 45.040 ;
        RECT 103.825 44.640 104.225 45.040 ;
        RECT 105.825 44.640 106.225 45.040 ;
        RECT 107.825 44.640 108.225 45.040 ;
        RECT 109.825 44.640 110.225 45.040 ;
        RECT 111.825 44.640 112.225 45.040 ;
        RECT 113.825 44.640 114.225 45.040 ;
        RECT 115.825 44.640 116.225 45.040 ;
        RECT 117.825 44.640 118.225 45.040 ;
        RECT 119.825 44.640 120.225 45.040 ;
        RECT 121.825 44.640 122.225 45.040 ;
        RECT 123.825 44.640 124.225 45.040 ;
        RECT 125.825 44.640 126.225 45.040 ;
        RECT 127.825 44.640 128.225 45.040 ;
        RECT 129.825 44.640 130.225 45.040 ;
        RECT 131.825 44.640 132.225 45.040 ;
        RECT 133.825 44.640 134.225 45.040 ;
        RECT 135.825 44.640 136.225 45.040 ;
        RECT 137.825 44.640 138.225 45.040 ;
        RECT 139.825 44.640 140.225 45.040 ;
        RECT 141.825 44.640 142.225 45.040 ;
        RECT 143.825 44.640 144.225 45.040 ;
        RECT 145.825 44.640 146.225 45.040 ;
        RECT 147.825 44.640 148.225 45.040 ;
        RECT 149.825 44.640 150.225 45.040 ;
        RECT 151.825 44.640 152.225 45.040 ;
        RECT 153.825 44.640 154.225 45.040 ;
        RECT 6.890 44.440 8.540 44.640 ;
        RECT 8.890 44.440 24.540 44.640 ;
        RECT 24.890 44.440 38.540 44.640 ;
        RECT 38.890 44.440 74.540 44.640 ;
        RECT 86.575 44.440 122.225 44.640 ;
        RECT 122.575 44.440 136.225 44.640 ;
        RECT 136.575 44.440 152.225 44.640 ;
        RECT 152.575 44.440 154.225 44.640 ;
        RECT 6.890 44.040 7.290 44.440 ;
        RECT 8.890 44.040 9.290 44.440 ;
        RECT 10.890 44.040 11.290 44.440 ;
        RECT 12.890 44.040 13.290 44.440 ;
        RECT 14.890 44.040 15.290 44.440 ;
        RECT 16.890 44.040 17.290 44.440 ;
        RECT 18.890 44.040 19.290 44.440 ;
        RECT 20.890 44.040 21.290 44.440 ;
        RECT 22.890 44.040 23.290 44.440 ;
        RECT 24.890 44.040 25.290 44.440 ;
        RECT 26.890 44.040 27.290 44.440 ;
        RECT 28.890 44.040 29.290 44.440 ;
        RECT 30.890 44.040 31.290 44.440 ;
        RECT 32.890 44.040 33.290 44.440 ;
        RECT 34.890 44.040 35.290 44.440 ;
        RECT 36.890 44.040 37.290 44.440 ;
        RECT 38.890 44.040 39.290 44.440 ;
        RECT 40.890 44.040 41.290 44.440 ;
        RECT 42.890 44.040 43.290 44.440 ;
        RECT 44.890 44.040 45.290 44.440 ;
        RECT 46.890 44.040 47.290 44.440 ;
        RECT 48.890 44.040 49.290 44.440 ;
        RECT 50.890 44.040 51.290 44.440 ;
        RECT 52.890 44.040 53.290 44.440 ;
        RECT 54.890 44.040 55.290 44.440 ;
        RECT 56.890 44.040 57.290 44.440 ;
        RECT 58.890 44.040 59.290 44.440 ;
        RECT 60.890 44.040 61.290 44.440 ;
        RECT 62.890 44.040 63.290 44.440 ;
        RECT 64.890 44.040 65.290 44.440 ;
        RECT 66.890 44.040 67.290 44.440 ;
        RECT 68.890 44.040 69.290 44.440 ;
        RECT 70.890 44.040 71.290 44.440 ;
        RECT 72.890 44.040 73.290 44.440 ;
        RECT 87.825 44.040 88.225 44.440 ;
        RECT 89.825 44.040 90.225 44.440 ;
        RECT 91.825 44.040 92.225 44.440 ;
        RECT 93.825 44.040 94.225 44.440 ;
        RECT 95.825 44.040 96.225 44.440 ;
        RECT 97.825 44.040 98.225 44.440 ;
        RECT 99.825 44.040 100.225 44.440 ;
        RECT 101.825 44.040 102.225 44.440 ;
        RECT 103.825 44.040 104.225 44.440 ;
        RECT 105.825 44.040 106.225 44.440 ;
        RECT 107.825 44.040 108.225 44.440 ;
        RECT 109.825 44.040 110.225 44.440 ;
        RECT 111.825 44.040 112.225 44.440 ;
        RECT 113.825 44.040 114.225 44.440 ;
        RECT 115.825 44.040 116.225 44.440 ;
        RECT 117.825 44.040 118.225 44.440 ;
        RECT 119.825 44.040 120.225 44.440 ;
        RECT 121.825 44.040 122.225 44.440 ;
        RECT 123.825 44.040 124.225 44.440 ;
        RECT 125.825 44.040 126.225 44.440 ;
        RECT 127.825 44.040 128.225 44.440 ;
        RECT 129.825 44.040 130.225 44.440 ;
        RECT 131.825 44.040 132.225 44.440 ;
        RECT 133.825 44.040 134.225 44.440 ;
        RECT 135.825 44.040 136.225 44.440 ;
        RECT 137.825 44.040 138.225 44.440 ;
        RECT 139.825 44.040 140.225 44.440 ;
        RECT 141.825 44.040 142.225 44.440 ;
        RECT 143.825 44.040 144.225 44.440 ;
        RECT 145.825 44.040 146.225 44.440 ;
        RECT 147.825 44.040 148.225 44.440 ;
        RECT 149.825 44.040 150.225 44.440 ;
        RECT 151.825 44.040 152.225 44.440 ;
        RECT 153.825 44.040 154.225 44.440 ;
        RECT 6.960 43.190 7.220 44.040 ;
        RECT 8.990 43.190 9.190 44.040 ;
        RECT 10.990 43.190 11.190 44.040 ;
        RECT 12.990 43.190 13.190 44.040 ;
        RECT 14.990 43.190 15.190 44.040 ;
        RECT 16.990 43.190 17.190 44.040 ;
        RECT 18.990 43.190 19.190 44.040 ;
        RECT 20.990 43.190 21.190 44.040 ;
        RECT 22.990 43.190 23.190 44.040 ;
        RECT 24.990 43.190 25.190 44.040 ;
        RECT 26.990 43.190 27.190 44.040 ;
        RECT 28.990 43.190 29.190 44.040 ;
        RECT 30.990 43.190 31.190 44.040 ;
        RECT 32.990 43.190 33.190 44.040 ;
        RECT 34.990 43.190 35.190 44.040 ;
        RECT 36.990 43.190 37.190 44.040 ;
        RECT 38.990 43.190 39.190 44.040 ;
        RECT 40.990 43.190 41.190 44.040 ;
        RECT 42.990 43.190 43.190 44.040 ;
        RECT 44.990 43.190 45.190 44.040 ;
        RECT 46.990 43.190 47.190 44.040 ;
        RECT 48.990 43.190 49.190 44.040 ;
        RECT 50.990 43.190 51.190 44.040 ;
        RECT 52.990 43.190 53.190 44.040 ;
        RECT 54.990 43.190 55.190 44.040 ;
        RECT 56.990 43.190 57.190 44.040 ;
        RECT 58.990 43.190 59.190 44.040 ;
        RECT 60.990 43.190 61.190 44.040 ;
        RECT 62.990 43.190 63.190 44.040 ;
        RECT 64.990 43.190 65.190 44.040 ;
        RECT 66.990 43.190 67.190 44.040 ;
        RECT 68.990 43.190 69.190 44.040 ;
        RECT 70.990 43.190 71.190 44.040 ;
        RECT 89.925 43.190 90.125 44.040 ;
        RECT 91.925 43.190 92.125 44.040 ;
        RECT 93.925 43.190 94.125 44.040 ;
        RECT 95.925 43.190 96.125 44.040 ;
        RECT 97.925 43.190 98.125 44.040 ;
        RECT 99.925 43.190 100.125 44.040 ;
        RECT 101.925 43.190 102.125 44.040 ;
        RECT 103.925 43.190 104.125 44.040 ;
        RECT 105.925 43.190 106.125 44.040 ;
        RECT 107.925 43.190 108.125 44.040 ;
        RECT 109.925 43.190 110.125 44.040 ;
        RECT 111.925 43.190 112.125 44.040 ;
        RECT 113.925 43.190 114.125 44.040 ;
        RECT 115.925 43.190 116.125 44.040 ;
        RECT 117.925 43.190 118.125 44.040 ;
        RECT 119.925 43.190 120.125 44.040 ;
        RECT 121.925 43.190 122.125 44.040 ;
        RECT 123.925 43.190 124.125 44.040 ;
        RECT 125.925 43.190 126.125 44.040 ;
        RECT 127.925 43.190 128.125 44.040 ;
        RECT 129.925 43.190 130.125 44.040 ;
        RECT 131.925 43.190 132.125 44.040 ;
        RECT 133.925 43.190 134.125 44.040 ;
        RECT 135.925 43.190 136.125 44.040 ;
        RECT 137.925 43.190 138.125 44.040 ;
        RECT 139.925 43.190 140.125 44.040 ;
        RECT 141.925 43.190 142.125 44.040 ;
        RECT 143.925 43.190 144.125 44.040 ;
        RECT 145.925 43.190 146.125 44.040 ;
        RECT 147.925 43.190 148.125 44.040 ;
        RECT 149.925 43.190 150.125 44.040 ;
        RECT 151.925 43.190 152.125 44.040 ;
        RECT 153.895 43.190 154.155 44.040 ;
        RECT 6.890 42.790 7.290 43.190 ;
        RECT 8.890 42.790 9.290 43.190 ;
        RECT 10.890 42.790 11.290 43.190 ;
        RECT 12.890 42.790 13.290 43.190 ;
        RECT 14.890 42.790 15.290 43.190 ;
        RECT 16.890 42.790 17.290 43.190 ;
        RECT 18.890 42.790 19.290 43.190 ;
        RECT 20.890 42.790 21.290 43.190 ;
        RECT 22.890 42.790 23.290 43.190 ;
        RECT 24.890 42.790 25.290 43.190 ;
        RECT 26.890 42.790 27.290 43.190 ;
        RECT 28.890 42.790 29.290 43.190 ;
        RECT 30.890 42.790 31.290 43.190 ;
        RECT 32.890 42.790 33.290 43.190 ;
        RECT 34.890 42.790 35.290 43.190 ;
        RECT 36.890 42.790 37.290 43.190 ;
        RECT 38.890 42.790 39.290 43.190 ;
        RECT 40.890 42.790 41.290 43.190 ;
        RECT 42.890 42.790 43.290 43.190 ;
        RECT 44.890 42.790 45.290 43.190 ;
        RECT 46.890 42.790 47.290 43.190 ;
        RECT 48.890 42.790 49.290 43.190 ;
        RECT 50.890 42.790 51.290 43.190 ;
        RECT 52.890 42.790 53.290 43.190 ;
        RECT 54.890 42.790 55.290 43.190 ;
        RECT 56.890 42.790 57.290 43.190 ;
        RECT 58.890 42.790 59.290 43.190 ;
        RECT 60.890 42.790 61.290 43.190 ;
        RECT 62.890 42.790 63.290 43.190 ;
        RECT 64.890 42.790 65.290 43.190 ;
        RECT 66.890 42.790 67.290 43.190 ;
        RECT 68.890 42.790 69.290 43.190 ;
        RECT 70.890 42.790 71.290 43.190 ;
        RECT 72.890 42.790 73.290 43.190 ;
        RECT 87.825 42.790 88.225 43.190 ;
        RECT 89.825 42.790 90.225 43.190 ;
        RECT 91.825 42.790 92.225 43.190 ;
        RECT 93.825 42.790 94.225 43.190 ;
        RECT 95.825 42.790 96.225 43.190 ;
        RECT 97.825 42.790 98.225 43.190 ;
        RECT 99.825 42.790 100.225 43.190 ;
        RECT 101.825 42.790 102.225 43.190 ;
        RECT 103.825 42.790 104.225 43.190 ;
        RECT 105.825 42.790 106.225 43.190 ;
        RECT 107.825 42.790 108.225 43.190 ;
        RECT 109.825 42.790 110.225 43.190 ;
        RECT 111.825 42.790 112.225 43.190 ;
        RECT 113.825 42.790 114.225 43.190 ;
        RECT 115.825 42.790 116.225 43.190 ;
        RECT 117.825 42.790 118.225 43.190 ;
        RECT 119.825 42.790 120.225 43.190 ;
        RECT 121.825 42.790 122.225 43.190 ;
        RECT 123.825 42.790 124.225 43.190 ;
        RECT 125.825 42.790 126.225 43.190 ;
        RECT 127.825 42.790 128.225 43.190 ;
        RECT 129.825 42.790 130.225 43.190 ;
        RECT 131.825 42.790 132.225 43.190 ;
        RECT 133.825 42.790 134.225 43.190 ;
        RECT 135.825 42.790 136.225 43.190 ;
        RECT 137.825 42.790 138.225 43.190 ;
        RECT 139.825 42.790 140.225 43.190 ;
        RECT 141.825 42.790 142.225 43.190 ;
        RECT 143.825 42.790 144.225 43.190 ;
        RECT 145.825 42.790 146.225 43.190 ;
        RECT 147.825 42.790 148.225 43.190 ;
        RECT 149.825 42.790 150.225 43.190 ;
        RECT 151.825 42.790 152.225 43.190 ;
        RECT 153.825 42.790 154.225 43.190 ;
        RECT 6.890 42.590 8.540 42.790 ;
        RECT 8.890 42.590 24.540 42.790 ;
        RECT 24.890 42.590 38.540 42.790 ;
        RECT 38.890 42.590 74.540 42.790 ;
        RECT 86.575 42.590 122.225 42.790 ;
        RECT 122.575 42.590 136.225 42.790 ;
        RECT 136.575 42.590 152.225 42.790 ;
        RECT 152.575 42.590 154.225 42.790 ;
        RECT 6.890 42.190 7.290 42.590 ;
        RECT 8.890 42.190 9.290 42.590 ;
        RECT 10.890 42.190 11.290 42.590 ;
        RECT 12.890 42.190 13.290 42.590 ;
        RECT 14.890 42.190 15.290 42.590 ;
        RECT 16.890 42.190 17.290 42.590 ;
        RECT 18.890 42.190 19.290 42.590 ;
        RECT 20.890 42.190 21.290 42.590 ;
        RECT 22.890 42.190 23.290 42.590 ;
        RECT 24.890 42.190 25.290 42.590 ;
        RECT 26.890 42.190 27.290 42.590 ;
        RECT 28.890 42.190 29.290 42.590 ;
        RECT 30.890 42.190 31.290 42.590 ;
        RECT 32.890 42.190 33.290 42.590 ;
        RECT 34.890 42.190 35.290 42.590 ;
        RECT 36.890 42.190 37.290 42.590 ;
        RECT 38.890 42.190 39.290 42.590 ;
        RECT 40.890 42.190 41.290 42.590 ;
        RECT 42.890 42.190 43.290 42.590 ;
        RECT 44.890 42.190 45.290 42.590 ;
        RECT 46.890 42.190 47.290 42.590 ;
        RECT 48.890 42.190 49.290 42.590 ;
        RECT 50.890 42.190 51.290 42.590 ;
        RECT 52.890 42.190 53.290 42.590 ;
        RECT 54.890 42.190 55.290 42.590 ;
        RECT 56.890 42.190 57.290 42.590 ;
        RECT 58.890 42.190 59.290 42.590 ;
        RECT 60.890 42.190 61.290 42.590 ;
        RECT 62.890 42.190 63.290 42.590 ;
        RECT 64.890 42.190 65.290 42.590 ;
        RECT 66.890 42.190 67.290 42.590 ;
        RECT 68.890 42.190 69.290 42.590 ;
        RECT 70.890 42.190 71.290 42.590 ;
        RECT 72.890 42.190 73.290 42.590 ;
        RECT 87.825 42.190 88.225 42.590 ;
        RECT 89.825 42.190 90.225 42.590 ;
        RECT 91.825 42.190 92.225 42.590 ;
        RECT 93.825 42.190 94.225 42.590 ;
        RECT 95.825 42.190 96.225 42.590 ;
        RECT 97.825 42.190 98.225 42.590 ;
        RECT 99.825 42.190 100.225 42.590 ;
        RECT 101.825 42.190 102.225 42.590 ;
        RECT 103.825 42.190 104.225 42.590 ;
        RECT 105.825 42.190 106.225 42.590 ;
        RECT 107.825 42.190 108.225 42.590 ;
        RECT 109.825 42.190 110.225 42.590 ;
        RECT 111.825 42.190 112.225 42.590 ;
        RECT 113.825 42.190 114.225 42.590 ;
        RECT 115.825 42.190 116.225 42.590 ;
        RECT 117.825 42.190 118.225 42.590 ;
        RECT 119.825 42.190 120.225 42.590 ;
        RECT 121.825 42.190 122.225 42.590 ;
        RECT 123.825 42.190 124.225 42.590 ;
        RECT 125.825 42.190 126.225 42.590 ;
        RECT 127.825 42.190 128.225 42.590 ;
        RECT 129.825 42.190 130.225 42.590 ;
        RECT 131.825 42.190 132.225 42.590 ;
        RECT 133.825 42.190 134.225 42.590 ;
        RECT 135.825 42.190 136.225 42.590 ;
        RECT 137.825 42.190 138.225 42.590 ;
        RECT 139.825 42.190 140.225 42.590 ;
        RECT 141.825 42.190 142.225 42.590 ;
        RECT 143.825 42.190 144.225 42.590 ;
        RECT 145.825 42.190 146.225 42.590 ;
        RECT 147.825 42.190 148.225 42.590 ;
        RECT 149.825 42.190 150.225 42.590 ;
        RECT 151.825 42.190 152.225 42.590 ;
        RECT 153.825 42.190 154.225 42.590 ;
        RECT 6.960 41.340 7.220 42.190 ;
        RECT 8.990 41.340 9.190 42.190 ;
        RECT 10.990 41.340 11.190 42.190 ;
        RECT 12.990 41.340 13.190 42.190 ;
        RECT 14.990 41.340 15.190 42.190 ;
        RECT 16.990 41.340 17.190 42.190 ;
        RECT 18.990 41.340 19.190 42.190 ;
        RECT 20.990 41.340 21.190 42.190 ;
        RECT 22.990 41.340 23.190 42.190 ;
        RECT 24.990 41.340 25.190 42.190 ;
        RECT 26.990 41.340 27.190 42.190 ;
        RECT 28.990 41.340 29.190 42.190 ;
        RECT 30.990 41.340 31.190 42.190 ;
        RECT 32.990 41.340 33.190 42.190 ;
        RECT 34.990 41.340 35.190 42.190 ;
        RECT 36.990 41.340 37.190 42.190 ;
        RECT 38.990 41.340 39.190 42.190 ;
        RECT 40.990 41.340 41.190 42.190 ;
        RECT 42.990 41.340 43.190 42.190 ;
        RECT 44.990 41.340 45.190 42.190 ;
        RECT 46.990 41.340 47.190 42.190 ;
        RECT 48.990 41.340 49.190 42.190 ;
        RECT 50.990 41.340 51.190 42.190 ;
        RECT 52.990 41.340 53.190 42.190 ;
        RECT 54.990 41.340 55.190 42.190 ;
        RECT 56.990 41.340 57.190 42.190 ;
        RECT 58.990 41.340 59.190 42.190 ;
        RECT 60.990 41.340 61.190 42.190 ;
        RECT 62.990 41.340 63.190 42.190 ;
        RECT 64.990 41.340 65.190 42.190 ;
        RECT 66.990 41.340 67.190 42.190 ;
        RECT 68.990 41.340 69.190 42.190 ;
        RECT 70.990 41.340 71.190 42.190 ;
        RECT 89.925 41.340 90.125 42.190 ;
        RECT 91.925 41.340 92.125 42.190 ;
        RECT 93.925 41.340 94.125 42.190 ;
        RECT 95.925 41.340 96.125 42.190 ;
        RECT 97.925 41.340 98.125 42.190 ;
        RECT 99.925 41.340 100.125 42.190 ;
        RECT 101.925 41.340 102.125 42.190 ;
        RECT 103.925 41.340 104.125 42.190 ;
        RECT 105.925 41.340 106.125 42.190 ;
        RECT 107.925 41.340 108.125 42.190 ;
        RECT 109.925 41.340 110.125 42.190 ;
        RECT 111.925 41.340 112.125 42.190 ;
        RECT 113.925 41.340 114.125 42.190 ;
        RECT 115.925 41.340 116.125 42.190 ;
        RECT 117.925 41.340 118.125 42.190 ;
        RECT 119.925 41.340 120.125 42.190 ;
        RECT 121.925 41.340 122.125 42.190 ;
        RECT 123.925 41.340 124.125 42.190 ;
        RECT 125.925 41.340 126.125 42.190 ;
        RECT 127.925 41.340 128.125 42.190 ;
        RECT 129.925 41.340 130.125 42.190 ;
        RECT 131.925 41.340 132.125 42.190 ;
        RECT 133.925 41.340 134.125 42.190 ;
        RECT 135.925 41.340 136.125 42.190 ;
        RECT 137.925 41.340 138.125 42.190 ;
        RECT 139.925 41.340 140.125 42.190 ;
        RECT 141.925 41.340 142.125 42.190 ;
        RECT 143.925 41.340 144.125 42.190 ;
        RECT 145.925 41.340 146.125 42.190 ;
        RECT 147.925 41.340 148.125 42.190 ;
        RECT 149.925 41.340 150.125 42.190 ;
        RECT 151.925 41.340 152.125 42.190 ;
        RECT 153.895 41.340 154.155 42.190 ;
        RECT 6.890 40.940 7.290 41.340 ;
        RECT 8.890 40.940 9.290 41.340 ;
        RECT 10.890 40.940 11.290 41.340 ;
        RECT 12.890 40.940 13.290 41.340 ;
        RECT 14.890 40.940 15.290 41.340 ;
        RECT 16.890 40.940 17.290 41.340 ;
        RECT 18.890 40.940 19.290 41.340 ;
        RECT 20.890 40.940 21.290 41.340 ;
        RECT 22.890 40.940 23.290 41.340 ;
        RECT 24.890 40.940 25.290 41.340 ;
        RECT 26.890 40.940 27.290 41.340 ;
        RECT 28.890 40.940 29.290 41.340 ;
        RECT 30.890 40.940 31.290 41.340 ;
        RECT 32.890 40.940 33.290 41.340 ;
        RECT 34.890 40.940 35.290 41.340 ;
        RECT 36.890 40.940 37.290 41.340 ;
        RECT 38.890 40.940 39.290 41.340 ;
        RECT 40.890 40.940 41.290 41.340 ;
        RECT 42.890 40.940 43.290 41.340 ;
        RECT 44.890 40.940 45.290 41.340 ;
        RECT 46.890 40.940 47.290 41.340 ;
        RECT 48.890 40.940 49.290 41.340 ;
        RECT 50.890 40.940 51.290 41.340 ;
        RECT 52.890 40.940 53.290 41.340 ;
        RECT 54.890 40.940 55.290 41.340 ;
        RECT 56.890 40.940 57.290 41.340 ;
        RECT 58.890 40.940 59.290 41.340 ;
        RECT 60.890 40.940 61.290 41.340 ;
        RECT 62.890 40.940 63.290 41.340 ;
        RECT 64.890 40.940 65.290 41.340 ;
        RECT 66.890 40.940 67.290 41.340 ;
        RECT 68.890 40.940 69.290 41.340 ;
        RECT 70.890 40.940 71.290 41.340 ;
        RECT 72.890 40.940 73.290 41.340 ;
        RECT 87.825 40.940 88.225 41.340 ;
        RECT 89.825 40.940 90.225 41.340 ;
        RECT 91.825 40.940 92.225 41.340 ;
        RECT 93.825 40.940 94.225 41.340 ;
        RECT 95.825 40.940 96.225 41.340 ;
        RECT 97.825 40.940 98.225 41.340 ;
        RECT 99.825 40.940 100.225 41.340 ;
        RECT 101.825 40.940 102.225 41.340 ;
        RECT 103.825 40.940 104.225 41.340 ;
        RECT 105.825 40.940 106.225 41.340 ;
        RECT 107.825 40.940 108.225 41.340 ;
        RECT 109.825 40.940 110.225 41.340 ;
        RECT 111.825 40.940 112.225 41.340 ;
        RECT 113.825 40.940 114.225 41.340 ;
        RECT 115.825 40.940 116.225 41.340 ;
        RECT 117.825 40.940 118.225 41.340 ;
        RECT 119.825 40.940 120.225 41.340 ;
        RECT 121.825 40.940 122.225 41.340 ;
        RECT 123.825 40.940 124.225 41.340 ;
        RECT 125.825 40.940 126.225 41.340 ;
        RECT 127.825 40.940 128.225 41.340 ;
        RECT 129.825 40.940 130.225 41.340 ;
        RECT 131.825 40.940 132.225 41.340 ;
        RECT 133.825 40.940 134.225 41.340 ;
        RECT 135.825 40.940 136.225 41.340 ;
        RECT 137.825 40.940 138.225 41.340 ;
        RECT 139.825 40.940 140.225 41.340 ;
        RECT 141.825 40.940 142.225 41.340 ;
        RECT 143.825 40.940 144.225 41.340 ;
        RECT 145.825 40.940 146.225 41.340 ;
        RECT 147.825 40.940 148.225 41.340 ;
        RECT 149.825 40.940 150.225 41.340 ;
        RECT 151.825 40.940 152.225 41.340 ;
        RECT 153.825 40.940 154.225 41.340 ;
        RECT 6.890 40.740 8.540 40.940 ;
        RECT 8.890 40.740 24.540 40.940 ;
        RECT 24.890 40.740 38.540 40.940 ;
        RECT 38.890 40.740 74.540 40.940 ;
        RECT 86.575 40.740 122.225 40.940 ;
        RECT 122.575 40.740 136.225 40.940 ;
        RECT 136.575 40.740 152.225 40.940 ;
        RECT 152.575 40.740 154.225 40.940 ;
        RECT 6.890 40.340 7.290 40.740 ;
        RECT 8.890 40.340 9.290 40.740 ;
        RECT 10.890 40.340 11.290 40.740 ;
        RECT 12.890 40.340 13.290 40.740 ;
        RECT 14.890 40.340 15.290 40.740 ;
        RECT 16.890 40.340 17.290 40.740 ;
        RECT 18.890 40.340 19.290 40.740 ;
        RECT 20.890 40.340 21.290 40.740 ;
        RECT 22.890 40.340 23.290 40.740 ;
        RECT 24.890 40.340 25.290 40.740 ;
        RECT 26.890 40.340 27.290 40.740 ;
        RECT 28.890 40.340 29.290 40.740 ;
        RECT 30.890 40.340 31.290 40.740 ;
        RECT 32.890 40.340 33.290 40.740 ;
        RECT 34.890 40.340 35.290 40.740 ;
        RECT 36.890 40.340 37.290 40.740 ;
        RECT 38.890 40.340 39.290 40.740 ;
        RECT 40.890 40.340 41.290 40.740 ;
        RECT 42.890 40.340 43.290 40.740 ;
        RECT 44.890 40.340 45.290 40.740 ;
        RECT 46.890 40.340 47.290 40.740 ;
        RECT 48.890 40.340 49.290 40.740 ;
        RECT 50.890 40.340 51.290 40.740 ;
        RECT 52.890 40.340 53.290 40.740 ;
        RECT 54.890 40.340 55.290 40.740 ;
        RECT 56.890 40.340 57.290 40.740 ;
        RECT 58.890 40.340 59.290 40.740 ;
        RECT 60.890 40.340 61.290 40.740 ;
        RECT 62.890 40.340 63.290 40.740 ;
        RECT 64.890 40.340 65.290 40.740 ;
        RECT 66.890 40.340 67.290 40.740 ;
        RECT 68.890 40.340 69.290 40.740 ;
        RECT 70.890 40.340 71.290 40.740 ;
        RECT 72.890 40.340 73.290 40.740 ;
        RECT 87.825 40.340 88.225 40.740 ;
        RECT 89.825 40.340 90.225 40.740 ;
        RECT 91.825 40.340 92.225 40.740 ;
        RECT 93.825 40.340 94.225 40.740 ;
        RECT 95.825 40.340 96.225 40.740 ;
        RECT 97.825 40.340 98.225 40.740 ;
        RECT 99.825 40.340 100.225 40.740 ;
        RECT 101.825 40.340 102.225 40.740 ;
        RECT 103.825 40.340 104.225 40.740 ;
        RECT 105.825 40.340 106.225 40.740 ;
        RECT 107.825 40.340 108.225 40.740 ;
        RECT 109.825 40.340 110.225 40.740 ;
        RECT 111.825 40.340 112.225 40.740 ;
        RECT 113.825 40.340 114.225 40.740 ;
        RECT 115.825 40.340 116.225 40.740 ;
        RECT 117.825 40.340 118.225 40.740 ;
        RECT 119.825 40.340 120.225 40.740 ;
        RECT 121.825 40.340 122.225 40.740 ;
        RECT 123.825 40.340 124.225 40.740 ;
        RECT 125.825 40.340 126.225 40.740 ;
        RECT 127.825 40.340 128.225 40.740 ;
        RECT 129.825 40.340 130.225 40.740 ;
        RECT 131.825 40.340 132.225 40.740 ;
        RECT 133.825 40.340 134.225 40.740 ;
        RECT 135.825 40.340 136.225 40.740 ;
        RECT 137.825 40.340 138.225 40.740 ;
        RECT 139.825 40.340 140.225 40.740 ;
        RECT 141.825 40.340 142.225 40.740 ;
        RECT 143.825 40.340 144.225 40.740 ;
        RECT 145.825 40.340 146.225 40.740 ;
        RECT 147.825 40.340 148.225 40.740 ;
        RECT 149.825 40.340 150.225 40.740 ;
        RECT 151.825 40.340 152.225 40.740 ;
        RECT 153.825 40.340 154.225 40.740 ;
        RECT 6.960 39.490 7.220 40.340 ;
        RECT 8.990 39.490 9.190 40.340 ;
        RECT 10.990 39.490 11.190 40.340 ;
        RECT 12.990 39.490 13.190 40.340 ;
        RECT 14.990 39.490 15.190 40.340 ;
        RECT 16.990 39.490 17.190 40.340 ;
        RECT 18.990 39.490 19.190 40.340 ;
        RECT 20.990 39.490 21.190 40.340 ;
        RECT 22.990 39.490 23.190 40.340 ;
        RECT 24.990 39.490 25.190 40.340 ;
        RECT 26.990 39.490 27.190 40.340 ;
        RECT 28.990 39.490 29.190 40.340 ;
        RECT 30.990 39.490 31.190 40.340 ;
        RECT 32.990 39.490 33.190 40.340 ;
        RECT 34.990 39.490 35.190 40.340 ;
        RECT 36.990 39.490 37.190 40.340 ;
        RECT 38.990 39.490 39.190 40.340 ;
        RECT 40.990 39.490 41.190 40.340 ;
        RECT 42.990 39.490 43.190 40.340 ;
        RECT 44.990 39.490 45.190 40.340 ;
        RECT 46.990 39.490 47.190 40.340 ;
        RECT 48.990 39.490 49.190 40.340 ;
        RECT 50.990 39.490 51.190 40.340 ;
        RECT 52.990 39.490 53.190 40.340 ;
        RECT 54.990 39.490 55.190 40.340 ;
        RECT 56.990 39.490 57.190 40.340 ;
        RECT 58.990 39.490 59.190 40.340 ;
        RECT 60.990 39.490 61.190 40.340 ;
        RECT 62.990 39.490 63.190 40.340 ;
        RECT 64.990 39.490 65.190 40.340 ;
        RECT 66.990 39.490 67.190 40.340 ;
        RECT 68.990 39.490 69.190 40.340 ;
        RECT 70.990 39.490 71.190 40.340 ;
        RECT 89.925 39.490 90.125 40.340 ;
        RECT 91.925 39.490 92.125 40.340 ;
        RECT 93.925 39.490 94.125 40.340 ;
        RECT 95.925 39.490 96.125 40.340 ;
        RECT 97.925 39.490 98.125 40.340 ;
        RECT 99.925 39.490 100.125 40.340 ;
        RECT 101.925 39.490 102.125 40.340 ;
        RECT 103.925 39.490 104.125 40.340 ;
        RECT 105.925 39.490 106.125 40.340 ;
        RECT 107.925 39.490 108.125 40.340 ;
        RECT 109.925 39.490 110.125 40.340 ;
        RECT 111.925 39.490 112.125 40.340 ;
        RECT 113.925 39.490 114.125 40.340 ;
        RECT 115.925 39.490 116.125 40.340 ;
        RECT 117.925 39.490 118.125 40.340 ;
        RECT 119.925 39.490 120.125 40.340 ;
        RECT 121.925 39.490 122.125 40.340 ;
        RECT 123.925 39.490 124.125 40.340 ;
        RECT 125.925 39.490 126.125 40.340 ;
        RECT 127.925 39.490 128.125 40.340 ;
        RECT 129.925 39.490 130.125 40.340 ;
        RECT 131.925 39.490 132.125 40.340 ;
        RECT 133.925 39.490 134.125 40.340 ;
        RECT 135.925 39.490 136.125 40.340 ;
        RECT 137.925 39.490 138.125 40.340 ;
        RECT 139.925 39.490 140.125 40.340 ;
        RECT 141.925 39.490 142.125 40.340 ;
        RECT 143.925 39.490 144.125 40.340 ;
        RECT 145.925 39.490 146.125 40.340 ;
        RECT 147.925 39.490 148.125 40.340 ;
        RECT 149.925 39.490 150.125 40.340 ;
        RECT 151.925 39.490 152.125 40.340 ;
        RECT 153.895 39.490 154.155 40.340 ;
        RECT 6.890 39.090 7.290 39.490 ;
        RECT 8.890 39.090 9.290 39.490 ;
        RECT 10.890 39.090 11.290 39.490 ;
        RECT 12.890 39.090 13.290 39.490 ;
        RECT 14.890 39.090 15.290 39.490 ;
        RECT 16.890 39.090 17.290 39.490 ;
        RECT 18.890 39.090 19.290 39.490 ;
        RECT 20.890 39.090 21.290 39.490 ;
        RECT 22.890 39.090 23.290 39.490 ;
        RECT 24.890 39.090 25.290 39.490 ;
        RECT 26.890 39.090 27.290 39.490 ;
        RECT 28.890 39.090 29.290 39.490 ;
        RECT 30.890 39.090 31.290 39.490 ;
        RECT 32.890 39.090 33.290 39.490 ;
        RECT 34.890 39.090 35.290 39.490 ;
        RECT 36.890 39.090 37.290 39.490 ;
        RECT 38.890 39.090 39.290 39.490 ;
        RECT 40.890 39.090 41.290 39.490 ;
        RECT 42.890 39.090 43.290 39.490 ;
        RECT 44.890 39.090 45.290 39.490 ;
        RECT 46.890 39.090 47.290 39.490 ;
        RECT 48.890 39.090 49.290 39.490 ;
        RECT 50.890 39.090 51.290 39.490 ;
        RECT 52.890 39.090 53.290 39.490 ;
        RECT 54.890 39.090 55.290 39.490 ;
        RECT 56.890 39.090 57.290 39.490 ;
        RECT 58.890 39.090 59.290 39.490 ;
        RECT 60.890 39.090 61.290 39.490 ;
        RECT 62.890 39.090 63.290 39.490 ;
        RECT 64.890 39.090 65.290 39.490 ;
        RECT 66.890 39.090 67.290 39.490 ;
        RECT 68.890 39.090 69.290 39.490 ;
        RECT 70.890 39.090 71.290 39.490 ;
        RECT 72.890 39.090 73.290 39.490 ;
        RECT 87.825 39.090 88.225 39.490 ;
        RECT 89.825 39.090 90.225 39.490 ;
        RECT 91.825 39.090 92.225 39.490 ;
        RECT 93.825 39.090 94.225 39.490 ;
        RECT 95.825 39.090 96.225 39.490 ;
        RECT 97.825 39.090 98.225 39.490 ;
        RECT 99.825 39.090 100.225 39.490 ;
        RECT 101.825 39.090 102.225 39.490 ;
        RECT 103.825 39.090 104.225 39.490 ;
        RECT 105.825 39.090 106.225 39.490 ;
        RECT 107.825 39.090 108.225 39.490 ;
        RECT 109.825 39.090 110.225 39.490 ;
        RECT 111.825 39.090 112.225 39.490 ;
        RECT 113.825 39.090 114.225 39.490 ;
        RECT 115.825 39.090 116.225 39.490 ;
        RECT 117.825 39.090 118.225 39.490 ;
        RECT 119.825 39.090 120.225 39.490 ;
        RECT 121.825 39.090 122.225 39.490 ;
        RECT 123.825 39.090 124.225 39.490 ;
        RECT 125.825 39.090 126.225 39.490 ;
        RECT 127.825 39.090 128.225 39.490 ;
        RECT 129.825 39.090 130.225 39.490 ;
        RECT 131.825 39.090 132.225 39.490 ;
        RECT 133.825 39.090 134.225 39.490 ;
        RECT 135.825 39.090 136.225 39.490 ;
        RECT 137.825 39.090 138.225 39.490 ;
        RECT 139.825 39.090 140.225 39.490 ;
        RECT 141.825 39.090 142.225 39.490 ;
        RECT 143.825 39.090 144.225 39.490 ;
        RECT 145.825 39.090 146.225 39.490 ;
        RECT 147.825 39.090 148.225 39.490 ;
        RECT 149.825 39.090 150.225 39.490 ;
        RECT 151.825 39.090 152.225 39.490 ;
        RECT 153.825 39.090 154.225 39.490 ;
        RECT 6.890 38.890 8.540 39.090 ;
        RECT 8.890 38.890 24.540 39.090 ;
        RECT 24.890 38.890 38.540 39.090 ;
        RECT 38.890 38.890 74.540 39.090 ;
        RECT 86.575 38.890 122.225 39.090 ;
        RECT 122.575 38.890 136.225 39.090 ;
        RECT 136.575 38.890 152.225 39.090 ;
        RECT 152.575 38.890 154.225 39.090 ;
        RECT 6.890 38.490 7.290 38.890 ;
        RECT 8.890 38.490 9.290 38.890 ;
        RECT 10.890 38.490 11.290 38.890 ;
        RECT 12.890 38.490 13.290 38.890 ;
        RECT 14.890 38.490 15.290 38.890 ;
        RECT 16.890 38.490 17.290 38.890 ;
        RECT 18.890 38.490 19.290 38.890 ;
        RECT 20.890 38.490 21.290 38.890 ;
        RECT 22.890 38.490 23.290 38.890 ;
        RECT 24.890 38.490 25.290 38.890 ;
        RECT 26.890 38.490 27.290 38.890 ;
        RECT 28.890 38.490 29.290 38.890 ;
        RECT 30.890 38.490 31.290 38.890 ;
        RECT 32.890 38.490 33.290 38.890 ;
        RECT 34.890 38.490 35.290 38.890 ;
        RECT 36.890 38.490 37.290 38.890 ;
        RECT 38.890 38.490 39.290 38.890 ;
        RECT 40.890 38.490 41.290 38.890 ;
        RECT 42.890 38.490 43.290 38.890 ;
        RECT 44.890 38.490 45.290 38.890 ;
        RECT 46.890 38.490 47.290 38.890 ;
        RECT 48.890 38.490 49.290 38.890 ;
        RECT 50.890 38.490 51.290 38.890 ;
        RECT 52.890 38.490 53.290 38.890 ;
        RECT 54.890 38.490 55.290 38.890 ;
        RECT 56.890 38.490 57.290 38.890 ;
        RECT 58.890 38.490 59.290 38.890 ;
        RECT 60.890 38.490 61.290 38.890 ;
        RECT 62.890 38.490 63.290 38.890 ;
        RECT 64.890 38.490 65.290 38.890 ;
        RECT 66.890 38.490 67.290 38.890 ;
        RECT 68.890 38.490 69.290 38.890 ;
        RECT 70.890 38.490 71.290 38.890 ;
        RECT 72.890 38.490 73.290 38.890 ;
        RECT 87.825 38.490 88.225 38.890 ;
        RECT 89.825 38.490 90.225 38.890 ;
        RECT 91.825 38.490 92.225 38.890 ;
        RECT 93.825 38.490 94.225 38.890 ;
        RECT 95.825 38.490 96.225 38.890 ;
        RECT 97.825 38.490 98.225 38.890 ;
        RECT 99.825 38.490 100.225 38.890 ;
        RECT 101.825 38.490 102.225 38.890 ;
        RECT 103.825 38.490 104.225 38.890 ;
        RECT 105.825 38.490 106.225 38.890 ;
        RECT 107.825 38.490 108.225 38.890 ;
        RECT 109.825 38.490 110.225 38.890 ;
        RECT 111.825 38.490 112.225 38.890 ;
        RECT 113.825 38.490 114.225 38.890 ;
        RECT 115.825 38.490 116.225 38.890 ;
        RECT 117.825 38.490 118.225 38.890 ;
        RECT 119.825 38.490 120.225 38.890 ;
        RECT 121.825 38.490 122.225 38.890 ;
        RECT 123.825 38.490 124.225 38.890 ;
        RECT 125.825 38.490 126.225 38.890 ;
        RECT 127.825 38.490 128.225 38.890 ;
        RECT 129.825 38.490 130.225 38.890 ;
        RECT 131.825 38.490 132.225 38.890 ;
        RECT 133.825 38.490 134.225 38.890 ;
        RECT 135.825 38.490 136.225 38.890 ;
        RECT 137.825 38.490 138.225 38.890 ;
        RECT 139.825 38.490 140.225 38.890 ;
        RECT 141.825 38.490 142.225 38.890 ;
        RECT 143.825 38.490 144.225 38.890 ;
        RECT 145.825 38.490 146.225 38.890 ;
        RECT 147.825 38.490 148.225 38.890 ;
        RECT 149.825 38.490 150.225 38.890 ;
        RECT 151.825 38.490 152.225 38.890 ;
        RECT 153.825 38.490 154.225 38.890 ;
        RECT 6.960 37.640 7.220 38.490 ;
        RECT 8.990 37.640 9.190 38.490 ;
        RECT 10.990 37.640 11.190 38.490 ;
        RECT 12.990 37.640 13.190 38.490 ;
        RECT 14.990 37.640 15.190 38.490 ;
        RECT 16.990 37.640 17.190 38.490 ;
        RECT 18.990 37.640 19.190 38.490 ;
        RECT 20.990 37.640 21.190 38.490 ;
        RECT 22.990 37.640 23.190 38.490 ;
        RECT 24.990 37.640 25.190 38.490 ;
        RECT 26.990 37.640 27.190 38.490 ;
        RECT 28.990 37.640 29.190 38.490 ;
        RECT 30.990 37.640 31.190 38.490 ;
        RECT 32.990 37.640 33.190 38.490 ;
        RECT 34.990 37.640 35.190 38.490 ;
        RECT 36.990 37.640 37.190 38.490 ;
        RECT 123.925 37.640 124.125 38.490 ;
        RECT 125.925 37.640 126.125 38.490 ;
        RECT 127.925 37.640 128.125 38.490 ;
        RECT 129.925 37.640 130.125 38.490 ;
        RECT 131.925 37.640 132.125 38.490 ;
        RECT 133.925 37.640 134.125 38.490 ;
        RECT 135.925 37.640 136.125 38.490 ;
        RECT 137.925 37.640 138.125 38.490 ;
        RECT 139.925 37.640 140.125 38.490 ;
        RECT 141.925 37.640 142.125 38.490 ;
        RECT 143.925 37.640 144.125 38.490 ;
        RECT 145.925 37.640 146.125 38.490 ;
        RECT 147.925 37.640 148.125 38.490 ;
        RECT 149.925 37.640 150.125 38.490 ;
        RECT 151.925 37.640 152.125 38.490 ;
        RECT 153.895 37.640 154.155 38.490 ;
        RECT 6.890 37.240 7.290 37.640 ;
        RECT 8.890 37.240 9.290 37.640 ;
        RECT 10.890 37.240 11.290 37.640 ;
        RECT 12.890 37.240 13.290 37.640 ;
        RECT 14.890 37.240 15.290 37.640 ;
        RECT 16.890 37.240 17.290 37.640 ;
        RECT 18.890 37.240 19.290 37.640 ;
        RECT 20.890 37.240 21.290 37.640 ;
        RECT 22.890 37.240 23.290 37.640 ;
        RECT 24.890 37.240 25.290 37.640 ;
        RECT 26.890 37.240 27.290 37.640 ;
        RECT 28.890 37.240 29.290 37.640 ;
        RECT 30.890 37.240 31.290 37.640 ;
        RECT 32.890 37.240 33.290 37.640 ;
        RECT 34.890 37.240 35.290 37.640 ;
        RECT 36.890 37.240 37.290 37.640 ;
        RECT 38.890 37.240 39.290 37.640 ;
        RECT 40.890 37.240 41.290 37.640 ;
        RECT 42.890 37.240 43.290 37.640 ;
        RECT 44.890 37.240 45.290 37.640 ;
        RECT 46.890 37.240 47.290 37.640 ;
        RECT 48.890 37.240 49.290 37.640 ;
        RECT 50.890 37.240 51.290 37.640 ;
        RECT 52.890 37.240 53.290 37.640 ;
        RECT 54.890 37.240 55.290 37.640 ;
        RECT 56.890 37.240 57.290 37.640 ;
        RECT 58.890 37.240 59.290 37.640 ;
        RECT 60.890 37.240 61.290 37.640 ;
        RECT 62.890 37.240 63.290 37.640 ;
        RECT 64.890 37.240 65.290 37.640 ;
        RECT 66.890 37.240 67.290 37.640 ;
        RECT 68.890 37.240 69.290 37.640 ;
        RECT 70.890 37.240 71.290 37.640 ;
        RECT 72.890 37.240 73.290 37.640 ;
        RECT 75.380 37.240 75.800 37.320 ;
        RECT 6.890 37.040 8.540 37.240 ;
        RECT 8.890 37.040 24.540 37.240 ;
        RECT 24.890 37.040 75.800 37.240 ;
        RECT 6.890 36.640 7.290 37.040 ;
        RECT 8.890 36.640 9.290 37.040 ;
        RECT 10.890 36.640 11.290 37.040 ;
        RECT 12.890 36.640 13.290 37.040 ;
        RECT 14.890 36.640 15.290 37.040 ;
        RECT 16.890 36.640 17.290 37.040 ;
        RECT 18.890 36.640 19.290 37.040 ;
        RECT 20.890 36.640 21.290 37.040 ;
        RECT 22.890 36.640 23.290 37.040 ;
        RECT 24.890 36.640 25.290 37.040 ;
        RECT 26.890 36.640 27.290 37.040 ;
        RECT 28.890 36.640 29.290 37.040 ;
        RECT 30.890 36.640 31.290 37.040 ;
        RECT 32.890 36.640 33.290 37.040 ;
        RECT 34.890 36.640 35.290 37.040 ;
        RECT 36.890 36.640 37.290 37.040 ;
        RECT 38.890 36.640 39.290 37.040 ;
        RECT 40.890 36.640 41.290 37.040 ;
        RECT 42.890 36.640 43.290 37.040 ;
        RECT 44.890 36.640 45.290 37.040 ;
        RECT 46.890 36.640 47.290 37.040 ;
        RECT 48.890 36.640 49.290 37.040 ;
        RECT 50.890 36.640 51.290 37.040 ;
        RECT 52.890 36.640 53.290 37.040 ;
        RECT 54.890 36.640 55.290 37.040 ;
        RECT 56.890 36.640 57.290 37.040 ;
        RECT 58.890 36.640 59.290 37.040 ;
        RECT 60.890 36.640 61.290 37.040 ;
        RECT 62.890 36.640 63.290 37.040 ;
        RECT 64.890 36.640 65.290 37.040 ;
        RECT 66.890 36.640 67.290 37.040 ;
        RECT 68.890 36.640 69.290 37.040 ;
        RECT 70.890 36.640 71.290 37.040 ;
        RECT 72.890 36.640 73.290 37.040 ;
        RECT 75.380 36.960 75.800 37.040 ;
        RECT 85.315 37.240 85.735 37.320 ;
        RECT 87.825 37.240 88.225 37.640 ;
        RECT 89.825 37.240 90.225 37.640 ;
        RECT 91.825 37.240 92.225 37.640 ;
        RECT 93.825 37.240 94.225 37.640 ;
        RECT 95.825 37.240 96.225 37.640 ;
        RECT 97.825 37.240 98.225 37.640 ;
        RECT 99.825 37.240 100.225 37.640 ;
        RECT 101.825 37.240 102.225 37.640 ;
        RECT 103.825 37.240 104.225 37.640 ;
        RECT 105.825 37.240 106.225 37.640 ;
        RECT 107.825 37.240 108.225 37.640 ;
        RECT 109.825 37.240 110.225 37.640 ;
        RECT 111.825 37.240 112.225 37.640 ;
        RECT 113.825 37.240 114.225 37.640 ;
        RECT 115.825 37.240 116.225 37.640 ;
        RECT 117.825 37.240 118.225 37.640 ;
        RECT 119.825 37.240 120.225 37.640 ;
        RECT 121.825 37.240 122.225 37.640 ;
        RECT 123.825 37.240 124.225 37.640 ;
        RECT 125.825 37.240 126.225 37.640 ;
        RECT 127.825 37.240 128.225 37.640 ;
        RECT 129.825 37.240 130.225 37.640 ;
        RECT 131.825 37.240 132.225 37.640 ;
        RECT 133.825 37.240 134.225 37.640 ;
        RECT 135.825 37.240 136.225 37.640 ;
        RECT 137.825 37.240 138.225 37.640 ;
        RECT 139.825 37.240 140.225 37.640 ;
        RECT 141.825 37.240 142.225 37.640 ;
        RECT 143.825 37.240 144.225 37.640 ;
        RECT 145.825 37.240 146.225 37.640 ;
        RECT 147.825 37.240 148.225 37.640 ;
        RECT 149.825 37.240 150.225 37.640 ;
        RECT 151.825 37.240 152.225 37.640 ;
        RECT 153.825 37.240 154.225 37.640 ;
        RECT 85.315 37.040 136.225 37.240 ;
        RECT 136.575 37.040 152.225 37.240 ;
        RECT 152.575 37.040 154.225 37.240 ;
        RECT 85.315 36.960 85.735 37.040 ;
        RECT 87.825 36.640 88.225 37.040 ;
        RECT 89.825 36.640 90.225 37.040 ;
        RECT 91.825 36.640 92.225 37.040 ;
        RECT 93.825 36.640 94.225 37.040 ;
        RECT 95.825 36.640 96.225 37.040 ;
        RECT 97.825 36.640 98.225 37.040 ;
        RECT 99.825 36.640 100.225 37.040 ;
        RECT 101.825 36.640 102.225 37.040 ;
        RECT 103.825 36.640 104.225 37.040 ;
        RECT 105.825 36.640 106.225 37.040 ;
        RECT 107.825 36.640 108.225 37.040 ;
        RECT 109.825 36.640 110.225 37.040 ;
        RECT 111.825 36.640 112.225 37.040 ;
        RECT 113.825 36.640 114.225 37.040 ;
        RECT 115.825 36.640 116.225 37.040 ;
        RECT 117.825 36.640 118.225 37.040 ;
        RECT 119.825 36.640 120.225 37.040 ;
        RECT 121.825 36.640 122.225 37.040 ;
        RECT 123.825 36.640 124.225 37.040 ;
        RECT 125.825 36.640 126.225 37.040 ;
        RECT 127.825 36.640 128.225 37.040 ;
        RECT 129.825 36.640 130.225 37.040 ;
        RECT 131.825 36.640 132.225 37.040 ;
        RECT 133.825 36.640 134.225 37.040 ;
        RECT 135.825 36.640 136.225 37.040 ;
        RECT 137.825 36.640 138.225 37.040 ;
        RECT 139.825 36.640 140.225 37.040 ;
        RECT 141.825 36.640 142.225 37.040 ;
        RECT 143.825 36.640 144.225 37.040 ;
        RECT 145.825 36.640 146.225 37.040 ;
        RECT 147.825 36.640 148.225 37.040 ;
        RECT 149.825 36.640 150.225 37.040 ;
        RECT 151.825 36.640 152.225 37.040 ;
        RECT 153.825 36.640 154.225 37.040 ;
        RECT 6.960 35.790 7.220 36.640 ;
        RECT 8.990 35.790 9.190 36.640 ;
        RECT 10.990 35.790 11.190 36.640 ;
        RECT 12.990 35.790 13.190 36.640 ;
        RECT 14.990 35.790 15.190 36.640 ;
        RECT 16.990 35.790 17.190 36.640 ;
        RECT 18.990 35.790 19.190 36.640 ;
        RECT 20.990 35.790 21.190 36.640 ;
        RECT 22.990 35.790 23.190 36.640 ;
        RECT 24.990 35.790 25.190 36.640 ;
        RECT 26.990 35.790 27.190 36.640 ;
        RECT 28.990 35.790 29.190 36.640 ;
        RECT 30.990 35.790 31.190 36.640 ;
        RECT 32.990 35.790 33.190 36.640 ;
        RECT 34.990 35.790 35.190 36.640 ;
        RECT 36.990 35.790 37.190 36.640 ;
        RECT 38.990 35.790 39.190 36.640 ;
        RECT 40.990 35.790 41.190 36.640 ;
        RECT 42.990 35.790 43.190 36.640 ;
        RECT 44.990 35.790 45.190 36.640 ;
        RECT 46.990 35.790 47.190 36.640 ;
        RECT 48.990 35.790 49.190 36.640 ;
        RECT 50.990 35.790 51.190 36.640 ;
        RECT 52.990 35.790 53.190 36.640 ;
        RECT 54.990 35.790 55.190 36.640 ;
        RECT 56.990 35.790 57.190 36.640 ;
        RECT 58.990 35.790 59.190 36.640 ;
        RECT 60.990 35.790 61.190 36.640 ;
        RECT 62.990 35.790 63.190 36.640 ;
        RECT 64.990 35.790 65.190 36.640 ;
        RECT 66.990 35.790 67.190 36.640 ;
        RECT 68.990 35.790 69.190 36.640 ;
        RECT 70.990 35.790 71.190 36.640 ;
        RECT 89.925 35.790 90.125 36.640 ;
        RECT 91.925 35.790 92.125 36.640 ;
        RECT 93.925 35.790 94.125 36.640 ;
        RECT 95.925 35.790 96.125 36.640 ;
        RECT 97.925 35.790 98.125 36.640 ;
        RECT 99.925 35.790 100.125 36.640 ;
        RECT 101.925 35.790 102.125 36.640 ;
        RECT 103.925 35.790 104.125 36.640 ;
        RECT 105.925 35.790 106.125 36.640 ;
        RECT 107.925 35.790 108.125 36.640 ;
        RECT 109.925 35.790 110.125 36.640 ;
        RECT 111.925 35.790 112.125 36.640 ;
        RECT 113.925 35.790 114.125 36.640 ;
        RECT 115.925 35.790 116.125 36.640 ;
        RECT 117.925 35.790 118.125 36.640 ;
        RECT 119.925 35.790 120.125 36.640 ;
        RECT 121.925 35.790 122.125 36.640 ;
        RECT 123.925 35.790 124.125 36.640 ;
        RECT 125.925 35.790 126.125 36.640 ;
        RECT 127.925 35.790 128.125 36.640 ;
        RECT 129.925 35.790 130.125 36.640 ;
        RECT 131.925 35.790 132.125 36.640 ;
        RECT 133.925 35.790 134.125 36.640 ;
        RECT 135.925 35.790 136.125 36.640 ;
        RECT 137.925 35.790 138.125 36.640 ;
        RECT 139.925 35.790 140.125 36.640 ;
        RECT 141.925 35.790 142.125 36.640 ;
        RECT 143.925 35.790 144.125 36.640 ;
        RECT 145.925 35.790 146.125 36.640 ;
        RECT 147.925 35.790 148.125 36.640 ;
        RECT 149.925 35.790 150.125 36.640 ;
        RECT 151.925 35.790 152.125 36.640 ;
        RECT 153.895 35.790 154.155 36.640 ;
        RECT 6.890 35.390 7.290 35.790 ;
        RECT 8.890 35.390 9.290 35.790 ;
        RECT 10.890 35.390 11.290 35.790 ;
        RECT 12.890 35.390 13.290 35.790 ;
        RECT 14.890 35.390 15.290 35.790 ;
        RECT 16.890 35.390 17.290 35.790 ;
        RECT 18.890 35.390 19.290 35.790 ;
        RECT 20.890 35.390 21.290 35.790 ;
        RECT 22.890 35.390 23.290 35.790 ;
        RECT 24.890 35.390 25.290 35.790 ;
        RECT 26.890 35.390 27.290 35.790 ;
        RECT 28.890 35.390 29.290 35.790 ;
        RECT 30.890 35.390 31.290 35.790 ;
        RECT 32.890 35.390 33.290 35.790 ;
        RECT 34.890 35.390 35.290 35.790 ;
        RECT 36.890 35.390 37.290 35.790 ;
        RECT 38.890 35.390 39.290 35.790 ;
        RECT 40.890 35.390 41.290 35.790 ;
        RECT 42.890 35.390 43.290 35.790 ;
        RECT 44.890 35.390 45.290 35.790 ;
        RECT 46.890 35.390 47.290 35.790 ;
        RECT 48.890 35.390 49.290 35.790 ;
        RECT 50.890 35.390 51.290 35.790 ;
        RECT 52.890 35.390 53.290 35.790 ;
        RECT 54.890 35.390 55.290 35.790 ;
        RECT 56.890 35.390 57.290 35.790 ;
        RECT 58.890 35.390 59.290 35.790 ;
        RECT 60.890 35.390 61.290 35.790 ;
        RECT 62.890 35.390 63.290 35.790 ;
        RECT 64.890 35.390 65.290 35.790 ;
        RECT 66.890 35.390 67.290 35.790 ;
        RECT 68.890 35.390 69.290 35.790 ;
        RECT 70.890 35.390 71.290 35.790 ;
        RECT 72.890 35.390 73.290 35.790 ;
        RECT 87.825 35.390 88.225 35.790 ;
        RECT 89.825 35.390 90.225 35.790 ;
        RECT 91.825 35.390 92.225 35.790 ;
        RECT 93.825 35.390 94.225 35.790 ;
        RECT 95.825 35.390 96.225 35.790 ;
        RECT 97.825 35.390 98.225 35.790 ;
        RECT 99.825 35.390 100.225 35.790 ;
        RECT 101.825 35.390 102.225 35.790 ;
        RECT 103.825 35.390 104.225 35.790 ;
        RECT 105.825 35.390 106.225 35.790 ;
        RECT 107.825 35.390 108.225 35.790 ;
        RECT 109.825 35.390 110.225 35.790 ;
        RECT 111.825 35.390 112.225 35.790 ;
        RECT 113.825 35.390 114.225 35.790 ;
        RECT 115.825 35.390 116.225 35.790 ;
        RECT 117.825 35.390 118.225 35.790 ;
        RECT 119.825 35.390 120.225 35.790 ;
        RECT 121.825 35.390 122.225 35.790 ;
        RECT 123.825 35.390 124.225 35.790 ;
        RECT 125.825 35.390 126.225 35.790 ;
        RECT 127.825 35.390 128.225 35.790 ;
        RECT 129.825 35.390 130.225 35.790 ;
        RECT 131.825 35.390 132.225 35.790 ;
        RECT 133.825 35.390 134.225 35.790 ;
        RECT 135.825 35.390 136.225 35.790 ;
        RECT 137.825 35.390 138.225 35.790 ;
        RECT 139.825 35.390 140.225 35.790 ;
        RECT 141.825 35.390 142.225 35.790 ;
        RECT 143.825 35.390 144.225 35.790 ;
        RECT 145.825 35.390 146.225 35.790 ;
        RECT 147.825 35.390 148.225 35.790 ;
        RECT 149.825 35.390 150.225 35.790 ;
        RECT 151.825 35.390 152.225 35.790 ;
        RECT 153.825 35.390 154.225 35.790 ;
        RECT 6.890 35.190 8.540 35.390 ;
        RECT 8.890 35.190 24.540 35.390 ;
        RECT 24.890 35.190 74.540 35.390 ;
        RECT 86.575 35.190 136.225 35.390 ;
        RECT 136.575 35.190 152.225 35.390 ;
        RECT 152.575 35.190 154.225 35.390 ;
        RECT 6.890 34.790 7.290 35.190 ;
        RECT 8.890 34.790 9.290 35.190 ;
        RECT 10.890 34.790 11.290 35.190 ;
        RECT 12.890 34.790 13.290 35.190 ;
        RECT 14.890 34.790 15.290 35.190 ;
        RECT 16.890 34.790 17.290 35.190 ;
        RECT 18.890 34.790 19.290 35.190 ;
        RECT 20.890 34.790 21.290 35.190 ;
        RECT 22.890 34.790 23.290 35.190 ;
        RECT 24.890 34.790 25.290 35.190 ;
        RECT 26.890 34.790 27.290 35.190 ;
        RECT 28.890 34.790 29.290 35.190 ;
        RECT 30.890 34.790 31.290 35.190 ;
        RECT 32.890 34.790 33.290 35.190 ;
        RECT 34.890 34.790 35.290 35.190 ;
        RECT 36.890 34.790 37.290 35.190 ;
        RECT 38.890 34.790 39.290 35.190 ;
        RECT 40.890 34.790 41.290 35.190 ;
        RECT 42.890 34.790 43.290 35.190 ;
        RECT 44.890 34.790 45.290 35.190 ;
        RECT 46.890 34.790 47.290 35.190 ;
        RECT 48.890 34.790 49.290 35.190 ;
        RECT 50.890 34.790 51.290 35.190 ;
        RECT 52.890 34.790 53.290 35.190 ;
        RECT 54.890 34.790 55.290 35.190 ;
        RECT 56.890 34.790 57.290 35.190 ;
        RECT 58.890 34.790 59.290 35.190 ;
        RECT 60.890 34.790 61.290 35.190 ;
        RECT 62.890 34.790 63.290 35.190 ;
        RECT 64.890 34.790 65.290 35.190 ;
        RECT 66.890 34.790 67.290 35.190 ;
        RECT 68.890 34.790 69.290 35.190 ;
        RECT 70.890 34.790 71.290 35.190 ;
        RECT 72.890 34.790 73.290 35.190 ;
        RECT 87.825 34.790 88.225 35.190 ;
        RECT 89.825 34.790 90.225 35.190 ;
        RECT 91.825 34.790 92.225 35.190 ;
        RECT 93.825 34.790 94.225 35.190 ;
        RECT 95.825 34.790 96.225 35.190 ;
        RECT 97.825 34.790 98.225 35.190 ;
        RECT 99.825 34.790 100.225 35.190 ;
        RECT 101.825 34.790 102.225 35.190 ;
        RECT 103.825 34.790 104.225 35.190 ;
        RECT 105.825 34.790 106.225 35.190 ;
        RECT 107.825 34.790 108.225 35.190 ;
        RECT 109.825 34.790 110.225 35.190 ;
        RECT 111.825 34.790 112.225 35.190 ;
        RECT 113.825 34.790 114.225 35.190 ;
        RECT 115.825 34.790 116.225 35.190 ;
        RECT 117.825 34.790 118.225 35.190 ;
        RECT 119.825 34.790 120.225 35.190 ;
        RECT 121.825 34.790 122.225 35.190 ;
        RECT 123.825 34.790 124.225 35.190 ;
        RECT 125.825 34.790 126.225 35.190 ;
        RECT 127.825 34.790 128.225 35.190 ;
        RECT 129.825 34.790 130.225 35.190 ;
        RECT 131.825 34.790 132.225 35.190 ;
        RECT 133.825 34.790 134.225 35.190 ;
        RECT 135.825 34.790 136.225 35.190 ;
        RECT 137.825 34.790 138.225 35.190 ;
        RECT 139.825 34.790 140.225 35.190 ;
        RECT 141.825 34.790 142.225 35.190 ;
        RECT 143.825 34.790 144.225 35.190 ;
        RECT 145.825 34.790 146.225 35.190 ;
        RECT 147.825 34.790 148.225 35.190 ;
        RECT 149.825 34.790 150.225 35.190 ;
        RECT 151.825 34.790 152.225 35.190 ;
        RECT 153.825 34.790 154.225 35.190 ;
        RECT 6.960 33.940 7.220 34.790 ;
        RECT 8.990 33.940 9.190 34.790 ;
        RECT 10.990 33.940 11.190 34.790 ;
        RECT 12.990 33.940 13.190 34.790 ;
        RECT 14.990 33.940 15.190 34.790 ;
        RECT 16.990 33.940 17.190 34.790 ;
        RECT 18.990 33.940 19.190 34.790 ;
        RECT 20.990 33.940 21.190 34.790 ;
        RECT 22.990 33.940 23.190 34.790 ;
        RECT 24.990 33.940 25.190 34.790 ;
        RECT 26.990 33.940 27.190 34.790 ;
        RECT 28.990 33.940 29.190 34.790 ;
        RECT 30.990 33.940 31.190 34.790 ;
        RECT 32.990 33.940 33.190 34.790 ;
        RECT 34.990 33.940 35.190 34.790 ;
        RECT 36.990 33.940 37.190 34.790 ;
        RECT 38.990 33.940 39.190 34.790 ;
        RECT 40.990 33.940 41.190 34.790 ;
        RECT 42.990 33.940 43.190 34.790 ;
        RECT 44.990 33.940 45.190 34.790 ;
        RECT 46.990 33.940 47.190 34.790 ;
        RECT 48.990 33.940 49.190 34.790 ;
        RECT 50.990 33.940 51.190 34.790 ;
        RECT 52.990 33.940 53.190 34.790 ;
        RECT 54.990 33.940 55.190 34.790 ;
        RECT 56.990 33.940 57.190 34.790 ;
        RECT 58.990 33.940 59.190 34.790 ;
        RECT 60.990 33.940 61.190 34.790 ;
        RECT 62.990 33.940 63.190 34.790 ;
        RECT 64.990 33.940 65.190 34.790 ;
        RECT 66.990 33.940 67.190 34.790 ;
        RECT 68.990 33.940 69.190 34.790 ;
        RECT 70.990 33.940 71.190 34.790 ;
        RECT 89.925 33.940 90.125 34.790 ;
        RECT 91.925 33.940 92.125 34.790 ;
        RECT 93.925 33.940 94.125 34.790 ;
        RECT 95.925 33.940 96.125 34.790 ;
        RECT 97.925 33.940 98.125 34.790 ;
        RECT 99.925 33.940 100.125 34.790 ;
        RECT 101.925 33.940 102.125 34.790 ;
        RECT 103.925 33.940 104.125 34.790 ;
        RECT 105.925 33.940 106.125 34.790 ;
        RECT 107.925 33.940 108.125 34.790 ;
        RECT 109.925 33.940 110.125 34.790 ;
        RECT 111.925 33.940 112.125 34.790 ;
        RECT 113.925 33.940 114.125 34.790 ;
        RECT 115.925 33.940 116.125 34.790 ;
        RECT 117.925 33.940 118.125 34.790 ;
        RECT 119.925 33.940 120.125 34.790 ;
        RECT 121.925 33.940 122.125 34.790 ;
        RECT 123.925 33.940 124.125 34.790 ;
        RECT 125.925 33.940 126.125 34.790 ;
        RECT 127.925 33.940 128.125 34.790 ;
        RECT 129.925 33.940 130.125 34.790 ;
        RECT 131.925 33.940 132.125 34.790 ;
        RECT 133.925 33.940 134.125 34.790 ;
        RECT 135.925 33.940 136.125 34.790 ;
        RECT 137.925 33.940 138.125 34.790 ;
        RECT 139.925 33.940 140.125 34.790 ;
        RECT 141.925 33.940 142.125 34.790 ;
        RECT 143.925 33.940 144.125 34.790 ;
        RECT 145.925 33.940 146.125 34.790 ;
        RECT 147.925 33.940 148.125 34.790 ;
        RECT 149.925 33.940 150.125 34.790 ;
        RECT 151.925 33.940 152.125 34.790 ;
        RECT 153.895 33.940 154.155 34.790 ;
        RECT 6.890 33.540 7.290 33.940 ;
        RECT 8.890 33.540 9.290 33.940 ;
        RECT 10.890 33.540 11.290 33.940 ;
        RECT 12.890 33.540 13.290 33.940 ;
        RECT 14.890 33.540 15.290 33.940 ;
        RECT 16.890 33.540 17.290 33.940 ;
        RECT 18.890 33.540 19.290 33.940 ;
        RECT 20.890 33.540 21.290 33.940 ;
        RECT 22.890 33.540 23.290 33.940 ;
        RECT 24.890 33.540 25.290 33.940 ;
        RECT 26.890 33.540 27.290 33.940 ;
        RECT 28.890 33.540 29.290 33.940 ;
        RECT 30.890 33.540 31.290 33.940 ;
        RECT 32.890 33.540 33.290 33.940 ;
        RECT 34.890 33.540 35.290 33.940 ;
        RECT 36.890 33.540 37.290 33.940 ;
        RECT 38.890 33.540 39.290 33.940 ;
        RECT 40.890 33.540 41.290 33.940 ;
        RECT 42.890 33.540 43.290 33.940 ;
        RECT 44.890 33.540 45.290 33.940 ;
        RECT 46.890 33.540 47.290 33.940 ;
        RECT 48.890 33.540 49.290 33.940 ;
        RECT 50.890 33.540 51.290 33.940 ;
        RECT 52.890 33.540 53.290 33.940 ;
        RECT 54.890 33.540 55.290 33.940 ;
        RECT 56.890 33.540 57.290 33.940 ;
        RECT 58.890 33.540 59.290 33.940 ;
        RECT 60.890 33.540 61.290 33.940 ;
        RECT 62.890 33.540 63.290 33.940 ;
        RECT 64.890 33.540 65.290 33.940 ;
        RECT 66.890 33.540 67.290 33.940 ;
        RECT 68.890 33.540 69.290 33.940 ;
        RECT 70.890 33.540 71.290 33.940 ;
        RECT 72.890 33.540 73.290 33.940 ;
        RECT 87.825 33.540 88.225 33.940 ;
        RECT 89.825 33.540 90.225 33.940 ;
        RECT 91.825 33.540 92.225 33.940 ;
        RECT 93.825 33.540 94.225 33.940 ;
        RECT 95.825 33.540 96.225 33.940 ;
        RECT 97.825 33.540 98.225 33.940 ;
        RECT 99.825 33.540 100.225 33.940 ;
        RECT 101.825 33.540 102.225 33.940 ;
        RECT 103.825 33.540 104.225 33.940 ;
        RECT 105.825 33.540 106.225 33.940 ;
        RECT 107.825 33.540 108.225 33.940 ;
        RECT 109.825 33.540 110.225 33.940 ;
        RECT 111.825 33.540 112.225 33.940 ;
        RECT 113.825 33.540 114.225 33.940 ;
        RECT 115.825 33.540 116.225 33.940 ;
        RECT 117.825 33.540 118.225 33.940 ;
        RECT 119.825 33.540 120.225 33.940 ;
        RECT 121.825 33.540 122.225 33.940 ;
        RECT 123.825 33.540 124.225 33.940 ;
        RECT 125.825 33.540 126.225 33.940 ;
        RECT 127.825 33.540 128.225 33.940 ;
        RECT 129.825 33.540 130.225 33.940 ;
        RECT 131.825 33.540 132.225 33.940 ;
        RECT 133.825 33.540 134.225 33.940 ;
        RECT 135.825 33.540 136.225 33.940 ;
        RECT 137.825 33.540 138.225 33.940 ;
        RECT 139.825 33.540 140.225 33.940 ;
        RECT 141.825 33.540 142.225 33.940 ;
        RECT 143.825 33.540 144.225 33.940 ;
        RECT 145.825 33.540 146.225 33.940 ;
        RECT 147.825 33.540 148.225 33.940 ;
        RECT 149.825 33.540 150.225 33.940 ;
        RECT 151.825 33.540 152.225 33.940 ;
        RECT 153.825 33.540 154.225 33.940 ;
        RECT 6.890 33.340 8.540 33.540 ;
        RECT 8.890 33.340 24.540 33.540 ;
        RECT 24.890 33.340 74.540 33.540 ;
        RECT 86.575 33.340 136.225 33.540 ;
        RECT 136.575 33.340 152.225 33.540 ;
        RECT 152.575 33.340 154.225 33.540 ;
        RECT 6.890 32.940 7.290 33.340 ;
        RECT 8.890 32.940 9.290 33.340 ;
        RECT 10.890 32.940 11.290 33.340 ;
        RECT 12.890 32.940 13.290 33.340 ;
        RECT 14.890 32.940 15.290 33.340 ;
        RECT 16.890 32.940 17.290 33.340 ;
        RECT 18.890 32.940 19.290 33.340 ;
        RECT 20.890 32.940 21.290 33.340 ;
        RECT 22.890 32.940 23.290 33.340 ;
        RECT 24.890 32.940 25.290 33.340 ;
        RECT 26.890 32.940 27.290 33.340 ;
        RECT 28.890 32.940 29.290 33.340 ;
        RECT 30.890 32.940 31.290 33.340 ;
        RECT 32.890 32.940 33.290 33.340 ;
        RECT 34.890 32.940 35.290 33.340 ;
        RECT 36.890 32.940 37.290 33.340 ;
        RECT 38.890 32.940 39.290 33.340 ;
        RECT 40.890 32.940 41.290 33.340 ;
        RECT 42.890 32.940 43.290 33.340 ;
        RECT 44.890 32.940 45.290 33.340 ;
        RECT 46.890 32.940 47.290 33.340 ;
        RECT 48.890 32.940 49.290 33.340 ;
        RECT 50.890 32.940 51.290 33.340 ;
        RECT 52.890 32.940 53.290 33.340 ;
        RECT 54.890 32.940 55.290 33.340 ;
        RECT 56.890 32.940 57.290 33.340 ;
        RECT 58.890 32.940 59.290 33.340 ;
        RECT 60.890 32.940 61.290 33.340 ;
        RECT 62.890 32.940 63.290 33.340 ;
        RECT 64.890 32.940 65.290 33.340 ;
        RECT 66.890 32.940 67.290 33.340 ;
        RECT 68.890 32.940 69.290 33.340 ;
        RECT 70.890 32.940 71.290 33.340 ;
        RECT 72.890 32.940 73.290 33.340 ;
        RECT 87.825 32.940 88.225 33.340 ;
        RECT 89.825 32.940 90.225 33.340 ;
        RECT 91.825 32.940 92.225 33.340 ;
        RECT 93.825 32.940 94.225 33.340 ;
        RECT 95.825 32.940 96.225 33.340 ;
        RECT 97.825 32.940 98.225 33.340 ;
        RECT 99.825 32.940 100.225 33.340 ;
        RECT 101.825 32.940 102.225 33.340 ;
        RECT 103.825 32.940 104.225 33.340 ;
        RECT 105.825 32.940 106.225 33.340 ;
        RECT 107.825 32.940 108.225 33.340 ;
        RECT 109.825 32.940 110.225 33.340 ;
        RECT 111.825 32.940 112.225 33.340 ;
        RECT 113.825 32.940 114.225 33.340 ;
        RECT 115.825 32.940 116.225 33.340 ;
        RECT 117.825 32.940 118.225 33.340 ;
        RECT 119.825 32.940 120.225 33.340 ;
        RECT 121.825 32.940 122.225 33.340 ;
        RECT 123.825 32.940 124.225 33.340 ;
        RECT 125.825 32.940 126.225 33.340 ;
        RECT 127.825 32.940 128.225 33.340 ;
        RECT 129.825 32.940 130.225 33.340 ;
        RECT 131.825 32.940 132.225 33.340 ;
        RECT 133.825 32.940 134.225 33.340 ;
        RECT 135.825 32.940 136.225 33.340 ;
        RECT 137.825 32.940 138.225 33.340 ;
        RECT 139.825 32.940 140.225 33.340 ;
        RECT 141.825 32.940 142.225 33.340 ;
        RECT 143.825 32.940 144.225 33.340 ;
        RECT 145.825 32.940 146.225 33.340 ;
        RECT 147.825 32.940 148.225 33.340 ;
        RECT 149.825 32.940 150.225 33.340 ;
        RECT 151.825 32.940 152.225 33.340 ;
        RECT 153.825 32.940 154.225 33.340 ;
        RECT 6.960 32.090 7.220 32.940 ;
        RECT 8.990 32.090 9.190 32.940 ;
        RECT 10.990 32.090 11.190 32.940 ;
        RECT 12.990 32.090 13.190 32.940 ;
        RECT 14.990 32.090 15.190 32.940 ;
        RECT 16.990 32.090 17.190 32.940 ;
        RECT 18.990 32.090 19.190 32.940 ;
        RECT 20.990 32.090 21.190 32.940 ;
        RECT 22.990 32.090 23.190 32.940 ;
        RECT 24.990 32.090 25.190 32.940 ;
        RECT 26.990 32.090 27.190 32.940 ;
        RECT 28.990 32.090 29.190 32.940 ;
        RECT 30.990 32.090 31.190 32.940 ;
        RECT 32.990 32.090 33.190 32.940 ;
        RECT 34.990 32.090 35.190 32.940 ;
        RECT 36.990 32.090 37.190 32.940 ;
        RECT 38.990 32.090 39.190 32.940 ;
        RECT 40.990 32.090 41.190 32.940 ;
        RECT 42.990 32.090 43.190 32.940 ;
        RECT 44.990 32.090 45.190 32.940 ;
        RECT 46.990 32.090 47.190 32.940 ;
        RECT 48.990 32.090 49.190 32.940 ;
        RECT 50.990 32.090 51.190 32.940 ;
        RECT 52.990 32.090 53.190 32.940 ;
        RECT 54.990 32.090 55.190 32.940 ;
        RECT 56.990 32.090 57.190 32.940 ;
        RECT 58.990 32.090 59.190 32.940 ;
        RECT 60.990 32.090 61.190 32.940 ;
        RECT 62.990 32.090 63.190 32.940 ;
        RECT 64.990 32.090 65.190 32.940 ;
        RECT 66.990 32.090 67.190 32.940 ;
        RECT 68.990 32.090 69.190 32.940 ;
        RECT 70.990 32.090 71.190 32.940 ;
        RECT 89.925 32.090 90.125 32.940 ;
        RECT 91.925 32.090 92.125 32.940 ;
        RECT 93.925 32.090 94.125 32.940 ;
        RECT 95.925 32.090 96.125 32.940 ;
        RECT 97.925 32.090 98.125 32.940 ;
        RECT 99.925 32.090 100.125 32.940 ;
        RECT 101.925 32.090 102.125 32.940 ;
        RECT 103.925 32.090 104.125 32.940 ;
        RECT 105.925 32.090 106.125 32.940 ;
        RECT 107.925 32.090 108.125 32.940 ;
        RECT 109.925 32.090 110.125 32.940 ;
        RECT 111.925 32.090 112.125 32.940 ;
        RECT 113.925 32.090 114.125 32.940 ;
        RECT 115.925 32.090 116.125 32.940 ;
        RECT 117.925 32.090 118.125 32.940 ;
        RECT 119.925 32.090 120.125 32.940 ;
        RECT 121.925 32.090 122.125 32.940 ;
        RECT 123.925 32.090 124.125 32.940 ;
        RECT 125.925 32.090 126.125 32.940 ;
        RECT 127.925 32.090 128.125 32.940 ;
        RECT 129.925 32.090 130.125 32.940 ;
        RECT 131.925 32.090 132.125 32.940 ;
        RECT 133.925 32.090 134.125 32.940 ;
        RECT 135.925 32.090 136.125 32.940 ;
        RECT 137.925 32.090 138.125 32.940 ;
        RECT 139.925 32.090 140.125 32.940 ;
        RECT 141.925 32.090 142.125 32.940 ;
        RECT 143.925 32.090 144.125 32.940 ;
        RECT 145.925 32.090 146.125 32.940 ;
        RECT 147.925 32.090 148.125 32.940 ;
        RECT 149.925 32.090 150.125 32.940 ;
        RECT 151.925 32.090 152.125 32.940 ;
        RECT 153.895 32.090 154.155 32.940 ;
        RECT 6.890 31.690 7.290 32.090 ;
        RECT 8.890 31.690 9.290 32.090 ;
        RECT 10.890 31.690 11.290 32.090 ;
        RECT 12.890 31.690 13.290 32.090 ;
        RECT 14.890 31.690 15.290 32.090 ;
        RECT 16.890 31.690 17.290 32.090 ;
        RECT 18.890 31.690 19.290 32.090 ;
        RECT 20.890 31.690 21.290 32.090 ;
        RECT 22.890 31.690 23.290 32.090 ;
        RECT 24.890 31.690 25.290 32.090 ;
        RECT 26.890 31.690 27.290 32.090 ;
        RECT 28.890 31.690 29.290 32.090 ;
        RECT 30.890 31.690 31.290 32.090 ;
        RECT 32.890 31.690 33.290 32.090 ;
        RECT 34.890 31.690 35.290 32.090 ;
        RECT 36.890 31.690 37.290 32.090 ;
        RECT 38.890 31.690 39.290 32.090 ;
        RECT 40.890 31.690 41.290 32.090 ;
        RECT 42.890 31.690 43.290 32.090 ;
        RECT 44.890 31.690 45.290 32.090 ;
        RECT 46.890 31.690 47.290 32.090 ;
        RECT 48.890 31.690 49.290 32.090 ;
        RECT 50.890 31.690 51.290 32.090 ;
        RECT 52.890 31.690 53.290 32.090 ;
        RECT 54.890 31.690 55.290 32.090 ;
        RECT 56.890 31.690 57.290 32.090 ;
        RECT 58.890 31.690 59.290 32.090 ;
        RECT 60.890 31.690 61.290 32.090 ;
        RECT 62.890 31.690 63.290 32.090 ;
        RECT 64.890 31.690 65.290 32.090 ;
        RECT 66.890 31.690 67.290 32.090 ;
        RECT 68.890 31.690 69.290 32.090 ;
        RECT 70.890 31.690 71.290 32.090 ;
        RECT 72.890 31.690 73.290 32.090 ;
        RECT 87.825 31.690 88.225 32.090 ;
        RECT 89.825 31.690 90.225 32.090 ;
        RECT 91.825 31.690 92.225 32.090 ;
        RECT 93.825 31.690 94.225 32.090 ;
        RECT 95.825 31.690 96.225 32.090 ;
        RECT 97.825 31.690 98.225 32.090 ;
        RECT 99.825 31.690 100.225 32.090 ;
        RECT 101.825 31.690 102.225 32.090 ;
        RECT 103.825 31.690 104.225 32.090 ;
        RECT 105.825 31.690 106.225 32.090 ;
        RECT 107.825 31.690 108.225 32.090 ;
        RECT 109.825 31.690 110.225 32.090 ;
        RECT 111.825 31.690 112.225 32.090 ;
        RECT 113.825 31.690 114.225 32.090 ;
        RECT 115.825 31.690 116.225 32.090 ;
        RECT 117.825 31.690 118.225 32.090 ;
        RECT 119.825 31.690 120.225 32.090 ;
        RECT 121.825 31.690 122.225 32.090 ;
        RECT 123.825 31.690 124.225 32.090 ;
        RECT 125.825 31.690 126.225 32.090 ;
        RECT 127.825 31.690 128.225 32.090 ;
        RECT 129.825 31.690 130.225 32.090 ;
        RECT 131.825 31.690 132.225 32.090 ;
        RECT 133.825 31.690 134.225 32.090 ;
        RECT 135.825 31.690 136.225 32.090 ;
        RECT 137.825 31.690 138.225 32.090 ;
        RECT 139.825 31.690 140.225 32.090 ;
        RECT 141.825 31.690 142.225 32.090 ;
        RECT 143.825 31.690 144.225 32.090 ;
        RECT 145.825 31.690 146.225 32.090 ;
        RECT 147.825 31.690 148.225 32.090 ;
        RECT 149.825 31.690 150.225 32.090 ;
        RECT 151.825 31.690 152.225 32.090 ;
        RECT 153.825 31.690 154.225 32.090 ;
        RECT 6.890 31.490 8.540 31.690 ;
        RECT 8.890 31.490 24.540 31.690 ;
        RECT 24.890 31.490 74.540 31.690 ;
        RECT 86.575 31.490 136.225 31.690 ;
        RECT 136.575 31.490 152.225 31.690 ;
        RECT 152.575 31.490 154.225 31.690 ;
        RECT 6.890 31.090 7.290 31.490 ;
        RECT 8.890 31.090 9.290 31.490 ;
        RECT 10.890 31.090 11.290 31.490 ;
        RECT 12.890 31.090 13.290 31.490 ;
        RECT 14.890 31.090 15.290 31.490 ;
        RECT 16.890 31.090 17.290 31.490 ;
        RECT 18.890 31.090 19.290 31.490 ;
        RECT 20.890 31.090 21.290 31.490 ;
        RECT 22.890 31.090 23.290 31.490 ;
        RECT 24.890 31.090 25.290 31.490 ;
        RECT 26.890 31.090 27.290 31.490 ;
        RECT 28.890 31.090 29.290 31.490 ;
        RECT 30.890 31.090 31.290 31.490 ;
        RECT 32.890 31.090 33.290 31.490 ;
        RECT 34.890 31.090 35.290 31.490 ;
        RECT 36.890 31.090 37.290 31.490 ;
        RECT 38.890 31.090 39.290 31.490 ;
        RECT 40.890 31.090 41.290 31.490 ;
        RECT 42.890 31.090 43.290 31.490 ;
        RECT 44.890 31.090 45.290 31.490 ;
        RECT 46.890 31.090 47.290 31.490 ;
        RECT 48.890 31.090 49.290 31.490 ;
        RECT 50.890 31.090 51.290 31.490 ;
        RECT 52.890 31.090 53.290 31.490 ;
        RECT 54.890 31.090 55.290 31.490 ;
        RECT 56.890 31.090 57.290 31.490 ;
        RECT 58.890 31.090 59.290 31.490 ;
        RECT 60.890 31.090 61.290 31.490 ;
        RECT 62.890 31.090 63.290 31.490 ;
        RECT 64.890 31.090 65.290 31.490 ;
        RECT 66.890 31.090 67.290 31.490 ;
        RECT 68.890 31.090 69.290 31.490 ;
        RECT 70.890 31.090 71.290 31.490 ;
        RECT 72.890 31.090 73.290 31.490 ;
        RECT 87.825 31.090 88.225 31.490 ;
        RECT 89.825 31.090 90.225 31.490 ;
        RECT 91.825 31.090 92.225 31.490 ;
        RECT 93.825 31.090 94.225 31.490 ;
        RECT 95.825 31.090 96.225 31.490 ;
        RECT 97.825 31.090 98.225 31.490 ;
        RECT 99.825 31.090 100.225 31.490 ;
        RECT 101.825 31.090 102.225 31.490 ;
        RECT 103.825 31.090 104.225 31.490 ;
        RECT 105.825 31.090 106.225 31.490 ;
        RECT 107.825 31.090 108.225 31.490 ;
        RECT 109.825 31.090 110.225 31.490 ;
        RECT 111.825 31.090 112.225 31.490 ;
        RECT 113.825 31.090 114.225 31.490 ;
        RECT 115.825 31.090 116.225 31.490 ;
        RECT 117.825 31.090 118.225 31.490 ;
        RECT 119.825 31.090 120.225 31.490 ;
        RECT 121.825 31.090 122.225 31.490 ;
        RECT 123.825 31.090 124.225 31.490 ;
        RECT 125.825 31.090 126.225 31.490 ;
        RECT 127.825 31.090 128.225 31.490 ;
        RECT 129.825 31.090 130.225 31.490 ;
        RECT 131.825 31.090 132.225 31.490 ;
        RECT 133.825 31.090 134.225 31.490 ;
        RECT 135.825 31.090 136.225 31.490 ;
        RECT 137.825 31.090 138.225 31.490 ;
        RECT 139.825 31.090 140.225 31.490 ;
        RECT 141.825 31.090 142.225 31.490 ;
        RECT 143.825 31.090 144.225 31.490 ;
        RECT 145.825 31.090 146.225 31.490 ;
        RECT 147.825 31.090 148.225 31.490 ;
        RECT 149.825 31.090 150.225 31.490 ;
        RECT 151.825 31.090 152.225 31.490 ;
        RECT 153.825 31.090 154.225 31.490 ;
        RECT 6.960 30.240 7.220 31.090 ;
        RECT 8.990 30.240 9.190 31.090 ;
        RECT 10.990 30.240 11.190 31.090 ;
        RECT 12.990 30.240 13.190 31.090 ;
        RECT 14.990 30.240 15.190 31.090 ;
        RECT 16.990 30.240 17.190 31.090 ;
        RECT 18.990 30.240 19.190 31.090 ;
        RECT 20.990 30.240 21.190 31.090 ;
        RECT 22.990 30.240 23.190 31.090 ;
        RECT 24.990 30.240 25.190 31.090 ;
        RECT 26.990 30.240 27.190 31.090 ;
        RECT 28.990 30.240 29.190 31.090 ;
        RECT 30.990 30.240 31.190 31.090 ;
        RECT 32.990 30.240 33.190 31.090 ;
        RECT 34.990 30.240 35.190 31.090 ;
        RECT 36.990 30.240 37.190 31.090 ;
        RECT 38.990 30.240 39.190 31.090 ;
        RECT 40.990 30.240 41.190 31.090 ;
        RECT 42.990 30.240 43.190 31.090 ;
        RECT 44.990 30.240 45.190 31.090 ;
        RECT 46.990 30.240 47.190 31.090 ;
        RECT 48.990 30.240 49.190 31.090 ;
        RECT 50.990 30.240 51.190 31.090 ;
        RECT 52.990 30.240 53.190 31.090 ;
        RECT 54.990 30.240 55.190 31.090 ;
        RECT 56.990 30.240 57.190 31.090 ;
        RECT 58.990 30.240 59.190 31.090 ;
        RECT 60.990 30.240 61.190 31.090 ;
        RECT 62.990 30.240 63.190 31.090 ;
        RECT 64.990 30.240 65.190 31.090 ;
        RECT 66.990 30.240 67.190 31.090 ;
        RECT 68.990 30.240 69.190 31.090 ;
        RECT 70.990 30.240 71.190 31.090 ;
        RECT 89.925 30.240 90.125 31.090 ;
        RECT 91.925 30.240 92.125 31.090 ;
        RECT 93.925 30.240 94.125 31.090 ;
        RECT 95.925 30.240 96.125 31.090 ;
        RECT 97.925 30.240 98.125 31.090 ;
        RECT 99.925 30.240 100.125 31.090 ;
        RECT 101.925 30.240 102.125 31.090 ;
        RECT 103.925 30.240 104.125 31.090 ;
        RECT 105.925 30.240 106.125 31.090 ;
        RECT 107.925 30.240 108.125 31.090 ;
        RECT 109.925 30.240 110.125 31.090 ;
        RECT 111.925 30.240 112.125 31.090 ;
        RECT 113.925 30.240 114.125 31.090 ;
        RECT 115.925 30.240 116.125 31.090 ;
        RECT 117.925 30.240 118.125 31.090 ;
        RECT 119.925 30.240 120.125 31.090 ;
        RECT 121.925 30.240 122.125 31.090 ;
        RECT 123.925 30.240 124.125 31.090 ;
        RECT 125.925 30.240 126.125 31.090 ;
        RECT 127.925 30.240 128.125 31.090 ;
        RECT 129.925 30.240 130.125 31.090 ;
        RECT 131.925 30.240 132.125 31.090 ;
        RECT 133.925 30.240 134.125 31.090 ;
        RECT 135.925 30.240 136.125 31.090 ;
        RECT 137.925 30.240 138.125 31.090 ;
        RECT 139.925 30.240 140.125 31.090 ;
        RECT 141.925 30.240 142.125 31.090 ;
        RECT 143.925 30.240 144.125 31.090 ;
        RECT 145.925 30.240 146.125 31.090 ;
        RECT 147.925 30.240 148.125 31.090 ;
        RECT 149.925 30.240 150.125 31.090 ;
        RECT 151.925 30.240 152.125 31.090 ;
        RECT 153.895 30.240 154.155 31.090 ;
        RECT 6.890 29.840 7.290 30.240 ;
        RECT 8.890 29.840 9.290 30.240 ;
        RECT 10.890 29.840 11.290 30.240 ;
        RECT 12.890 29.840 13.290 30.240 ;
        RECT 14.890 29.840 15.290 30.240 ;
        RECT 16.890 29.840 17.290 30.240 ;
        RECT 18.890 29.840 19.290 30.240 ;
        RECT 20.890 29.840 21.290 30.240 ;
        RECT 22.890 29.840 23.290 30.240 ;
        RECT 24.890 29.840 25.290 30.240 ;
        RECT 26.890 29.840 27.290 30.240 ;
        RECT 28.890 29.840 29.290 30.240 ;
        RECT 30.890 29.840 31.290 30.240 ;
        RECT 32.890 29.840 33.290 30.240 ;
        RECT 34.890 29.840 35.290 30.240 ;
        RECT 36.890 29.840 37.290 30.240 ;
        RECT 38.890 29.840 39.290 30.240 ;
        RECT 40.890 29.840 41.290 30.240 ;
        RECT 42.890 29.840 43.290 30.240 ;
        RECT 44.890 29.840 45.290 30.240 ;
        RECT 46.890 29.840 47.290 30.240 ;
        RECT 48.890 29.840 49.290 30.240 ;
        RECT 50.890 29.840 51.290 30.240 ;
        RECT 52.890 29.840 53.290 30.240 ;
        RECT 54.890 29.840 55.290 30.240 ;
        RECT 56.890 29.840 57.290 30.240 ;
        RECT 58.890 29.840 59.290 30.240 ;
        RECT 60.890 29.840 61.290 30.240 ;
        RECT 62.890 29.840 63.290 30.240 ;
        RECT 64.890 29.840 65.290 30.240 ;
        RECT 66.890 29.840 67.290 30.240 ;
        RECT 68.890 29.840 69.290 30.240 ;
        RECT 70.890 29.840 71.290 30.240 ;
        RECT 72.890 29.840 73.290 30.240 ;
        RECT 87.825 29.840 88.225 30.240 ;
        RECT 89.825 29.840 90.225 30.240 ;
        RECT 91.825 29.840 92.225 30.240 ;
        RECT 93.825 29.840 94.225 30.240 ;
        RECT 95.825 29.840 96.225 30.240 ;
        RECT 97.825 29.840 98.225 30.240 ;
        RECT 99.825 29.840 100.225 30.240 ;
        RECT 101.825 29.840 102.225 30.240 ;
        RECT 103.825 29.840 104.225 30.240 ;
        RECT 105.825 29.840 106.225 30.240 ;
        RECT 107.825 29.840 108.225 30.240 ;
        RECT 109.825 29.840 110.225 30.240 ;
        RECT 111.825 29.840 112.225 30.240 ;
        RECT 113.825 29.840 114.225 30.240 ;
        RECT 115.825 29.840 116.225 30.240 ;
        RECT 117.825 29.840 118.225 30.240 ;
        RECT 119.825 29.840 120.225 30.240 ;
        RECT 121.825 29.840 122.225 30.240 ;
        RECT 123.825 29.840 124.225 30.240 ;
        RECT 125.825 29.840 126.225 30.240 ;
        RECT 127.825 29.840 128.225 30.240 ;
        RECT 129.825 29.840 130.225 30.240 ;
        RECT 131.825 29.840 132.225 30.240 ;
        RECT 133.825 29.840 134.225 30.240 ;
        RECT 135.825 29.840 136.225 30.240 ;
        RECT 137.825 29.840 138.225 30.240 ;
        RECT 139.825 29.840 140.225 30.240 ;
        RECT 141.825 29.840 142.225 30.240 ;
        RECT 143.825 29.840 144.225 30.240 ;
        RECT 145.825 29.840 146.225 30.240 ;
        RECT 147.825 29.840 148.225 30.240 ;
        RECT 149.825 29.840 150.225 30.240 ;
        RECT 151.825 29.840 152.225 30.240 ;
        RECT 153.825 29.840 154.225 30.240 ;
        RECT 6.890 29.640 8.540 29.840 ;
        RECT 8.890 29.640 24.540 29.840 ;
        RECT 24.890 29.640 74.540 29.840 ;
        RECT 86.575 29.640 136.225 29.840 ;
        RECT 136.575 29.640 152.225 29.840 ;
        RECT 152.575 29.640 154.225 29.840 ;
        RECT 6.890 29.240 7.290 29.640 ;
        RECT 8.890 29.240 9.290 29.640 ;
        RECT 10.890 29.240 11.290 29.640 ;
        RECT 12.890 29.240 13.290 29.640 ;
        RECT 14.890 29.240 15.290 29.640 ;
        RECT 16.890 29.240 17.290 29.640 ;
        RECT 18.890 29.240 19.290 29.640 ;
        RECT 20.890 29.240 21.290 29.640 ;
        RECT 22.890 29.240 23.290 29.640 ;
        RECT 24.890 29.240 25.290 29.640 ;
        RECT 26.890 29.240 27.290 29.640 ;
        RECT 28.890 29.240 29.290 29.640 ;
        RECT 30.890 29.240 31.290 29.640 ;
        RECT 32.890 29.240 33.290 29.640 ;
        RECT 34.890 29.240 35.290 29.640 ;
        RECT 36.890 29.240 37.290 29.640 ;
        RECT 38.890 29.240 39.290 29.640 ;
        RECT 40.890 29.240 41.290 29.640 ;
        RECT 42.890 29.240 43.290 29.640 ;
        RECT 44.890 29.240 45.290 29.640 ;
        RECT 46.890 29.240 47.290 29.640 ;
        RECT 48.890 29.240 49.290 29.640 ;
        RECT 50.890 29.240 51.290 29.640 ;
        RECT 52.890 29.240 53.290 29.640 ;
        RECT 54.890 29.240 55.290 29.640 ;
        RECT 56.890 29.240 57.290 29.640 ;
        RECT 58.890 29.240 59.290 29.640 ;
        RECT 60.890 29.240 61.290 29.640 ;
        RECT 62.890 29.240 63.290 29.640 ;
        RECT 64.890 29.240 65.290 29.640 ;
        RECT 66.890 29.240 67.290 29.640 ;
        RECT 68.890 29.240 69.290 29.640 ;
        RECT 70.890 29.240 71.290 29.640 ;
        RECT 72.890 29.240 73.290 29.640 ;
        RECT 87.825 29.240 88.225 29.640 ;
        RECT 89.825 29.240 90.225 29.640 ;
        RECT 91.825 29.240 92.225 29.640 ;
        RECT 93.825 29.240 94.225 29.640 ;
        RECT 95.825 29.240 96.225 29.640 ;
        RECT 97.825 29.240 98.225 29.640 ;
        RECT 99.825 29.240 100.225 29.640 ;
        RECT 101.825 29.240 102.225 29.640 ;
        RECT 103.825 29.240 104.225 29.640 ;
        RECT 105.825 29.240 106.225 29.640 ;
        RECT 107.825 29.240 108.225 29.640 ;
        RECT 109.825 29.240 110.225 29.640 ;
        RECT 111.825 29.240 112.225 29.640 ;
        RECT 113.825 29.240 114.225 29.640 ;
        RECT 115.825 29.240 116.225 29.640 ;
        RECT 117.825 29.240 118.225 29.640 ;
        RECT 119.825 29.240 120.225 29.640 ;
        RECT 121.825 29.240 122.225 29.640 ;
        RECT 123.825 29.240 124.225 29.640 ;
        RECT 125.825 29.240 126.225 29.640 ;
        RECT 127.825 29.240 128.225 29.640 ;
        RECT 129.825 29.240 130.225 29.640 ;
        RECT 131.825 29.240 132.225 29.640 ;
        RECT 133.825 29.240 134.225 29.640 ;
        RECT 135.825 29.240 136.225 29.640 ;
        RECT 137.825 29.240 138.225 29.640 ;
        RECT 139.825 29.240 140.225 29.640 ;
        RECT 141.825 29.240 142.225 29.640 ;
        RECT 143.825 29.240 144.225 29.640 ;
        RECT 145.825 29.240 146.225 29.640 ;
        RECT 147.825 29.240 148.225 29.640 ;
        RECT 149.825 29.240 150.225 29.640 ;
        RECT 151.825 29.240 152.225 29.640 ;
        RECT 153.825 29.240 154.225 29.640 ;
        RECT 6.960 28.390 7.220 29.240 ;
        RECT 8.990 28.390 9.190 29.240 ;
        RECT 10.990 28.390 11.190 29.240 ;
        RECT 12.990 28.390 13.190 29.240 ;
        RECT 14.990 28.390 15.190 29.240 ;
        RECT 16.990 28.390 17.190 29.240 ;
        RECT 18.990 28.390 19.190 29.240 ;
        RECT 20.990 28.390 21.190 29.240 ;
        RECT 22.990 28.390 23.190 29.240 ;
        RECT 24.990 28.390 25.190 29.240 ;
        RECT 26.990 28.390 27.190 29.240 ;
        RECT 28.990 28.390 29.190 29.240 ;
        RECT 30.990 28.390 31.190 29.240 ;
        RECT 32.990 28.390 33.190 29.240 ;
        RECT 34.990 28.390 35.190 29.240 ;
        RECT 36.990 28.390 37.190 29.240 ;
        RECT 38.990 28.390 39.190 29.240 ;
        RECT 40.990 28.390 41.190 29.240 ;
        RECT 42.990 28.390 43.190 29.240 ;
        RECT 44.990 28.390 45.190 29.240 ;
        RECT 46.990 28.390 47.190 29.240 ;
        RECT 48.990 28.390 49.190 29.240 ;
        RECT 50.990 28.390 51.190 29.240 ;
        RECT 52.990 28.390 53.190 29.240 ;
        RECT 54.990 28.390 55.190 29.240 ;
        RECT 56.990 28.390 57.190 29.240 ;
        RECT 58.990 28.390 59.190 29.240 ;
        RECT 60.990 28.390 61.190 29.240 ;
        RECT 62.990 28.390 63.190 29.240 ;
        RECT 64.990 28.390 65.190 29.240 ;
        RECT 66.990 28.390 67.190 29.240 ;
        RECT 68.990 28.390 69.190 29.240 ;
        RECT 70.990 28.390 71.190 29.240 ;
        RECT 89.925 28.390 90.125 29.240 ;
        RECT 91.925 28.390 92.125 29.240 ;
        RECT 93.925 28.390 94.125 29.240 ;
        RECT 95.925 28.390 96.125 29.240 ;
        RECT 97.925 28.390 98.125 29.240 ;
        RECT 99.925 28.390 100.125 29.240 ;
        RECT 101.925 28.390 102.125 29.240 ;
        RECT 103.925 28.390 104.125 29.240 ;
        RECT 105.925 28.390 106.125 29.240 ;
        RECT 107.925 28.390 108.125 29.240 ;
        RECT 109.925 28.390 110.125 29.240 ;
        RECT 111.925 28.390 112.125 29.240 ;
        RECT 113.925 28.390 114.125 29.240 ;
        RECT 115.925 28.390 116.125 29.240 ;
        RECT 117.925 28.390 118.125 29.240 ;
        RECT 119.925 28.390 120.125 29.240 ;
        RECT 121.925 28.390 122.125 29.240 ;
        RECT 123.925 28.390 124.125 29.240 ;
        RECT 125.925 28.390 126.125 29.240 ;
        RECT 127.925 28.390 128.125 29.240 ;
        RECT 129.925 28.390 130.125 29.240 ;
        RECT 131.925 28.390 132.125 29.240 ;
        RECT 133.925 28.390 134.125 29.240 ;
        RECT 135.925 28.390 136.125 29.240 ;
        RECT 137.925 28.390 138.125 29.240 ;
        RECT 139.925 28.390 140.125 29.240 ;
        RECT 141.925 28.390 142.125 29.240 ;
        RECT 143.925 28.390 144.125 29.240 ;
        RECT 145.925 28.390 146.125 29.240 ;
        RECT 147.925 28.390 148.125 29.240 ;
        RECT 149.925 28.390 150.125 29.240 ;
        RECT 151.925 28.390 152.125 29.240 ;
        RECT 153.895 28.390 154.155 29.240 ;
        RECT 6.890 27.990 7.290 28.390 ;
        RECT 8.890 27.990 9.290 28.390 ;
        RECT 10.890 27.990 11.290 28.390 ;
        RECT 12.890 27.990 13.290 28.390 ;
        RECT 14.890 27.990 15.290 28.390 ;
        RECT 16.890 27.990 17.290 28.390 ;
        RECT 18.890 27.990 19.290 28.390 ;
        RECT 20.890 27.990 21.290 28.390 ;
        RECT 22.890 27.990 23.290 28.390 ;
        RECT 24.890 27.990 25.290 28.390 ;
        RECT 26.890 27.990 27.290 28.390 ;
        RECT 28.890 27.990 29.290 28.390 ;
        RECT 30.890 27.990 31.290 28.390 ;
        RECT 32.890 27.990 33.290 28.390 ;
        RECT 34.890 27.990 35.290 28.390 ;
        RECT 36.890 27.990 37.290 28.390 ;
        RECT 38.890 27.990 39.290 28.390 ;
        RECT 40.890 27.990 41.290 28.390 ;
        RECT 42.890 27.990 43.290 28.390 ;
        RECT 44.890 27.990 45.290 28.390 ;
        RECT 46.890 27.990 47.290 28.390 ;
        RECT 48.890 27.990 49.290 28.390 ;
        RECT 50.890 27.990 51.290 28.390 ;
        RECT 52.890 27.990 53.290 28.390 ;
        RECT 54.890 27.990 55.290 28.390 ;
        RECT 56.890 27.990 57.290 28.390 ;
        RECT 58.890 27.990 59.290 28.390 ;
        RECT 60.890 27.990 61.290 28.390 ;
        RECT 62.890 27.990 63.290 28.390 ;
        RECT 64.890 27.990 65.290 28.390 ;
        RECT 66.890 27.990 67.290 28.390 ;
        RECT 68.890 27.990 69.290 28.390 ;
        RECT 70.890 27.990 71.290 28.390 ;
        RECT 72.890 27.990 73.290 28.390 ;
        RECT 87.825 27.990 88.225 28.390 ;
        RECT 89.825 27.990 90.225 28.390 ;
        RECT 91.825 27.990 92.225 28.390 ;
        RECT 93.825 27.990 94.225 28.390 ;
        RECT 95.825 27.990 96.225 28.390 ;
        RECT 97.825 27.990 98.225 28.390 ;
        RECT 99.825 27.990 100.225 28.390 ;
        RECT 101.825 27.990 102.225 28.390 ;
        RECT 103.825 27.990 104.225 28.390 ;
        RECT 105.825 27.990 106.225 28.390 ;
        RECT 107.825 27.990 108.225 28.390 ;
        RECT 109.825 27.990 110.225 28.390 ;
        RECT 111.825 27.990 112.225 28.390 ;
        RECT 113.825 27.990 114.225 28.390 ;
        RECT 115.825 27.990 116.225 28.390 ;
        RECT 117.825 27.990 118.225 28.390 ;
        RECT 119.825 27.990 120.225 28.390 ;
        RECT 121.825 27.990 122.225 28.390 ;
        RECT 123.825 27.990 124.225 28.390 ;
        RECT 125.825 27.990 126.225 28.390 ;
        RECT 127.825 27.990 128.225 28.390 ;
        RECT 129.825 27.990 130.225 28.390 ;
        RECT 131.825 27.990 132.225 28.390 ;
        RECT 133.825 27.990 134.225 28.390 ;
        RECT 135.825 27.990 136.225 28.390 ;
        RECT 137.825 27.990 138.225 28.390 ;
        RECT 139.825 27.990 140.225 28.390 ;
        RECT 141.825 27.990 142.225 28.390 ;
        RECT 143.825 27.990 144.225 28.390 ;
        RECT 145.825 27.990 146.225 28.390 ;
        RECT 147.825 27.990 148.225 28.390 ;
        RECT 149.825 27.990 150.225 28.390 ;
        RECT 151.825 27.990 152.225 28.390 ;
        RECT 153.825 27.990 154.225 28.390 ;
        RECT 6.890 27.790 8.540 27.990 ;
        RECT 8.890 27.790 24.540 27.990 ;
        RECT 24.890 27.790 74.540 27.990 ;
        RECT 86.575 27.790 136.225 27.990 ;
        RECT 136.575 27.790 152.225 27.990 ;
        RECT 152.575 27.790 154.225 27.990 ;
        RECT 6.890 27.390 7.290 27.790 ;
        RECT 8.890 27.390 9.290 27.790 ;
        RECT 10.890 27.390 11.290 27.790 ;
        RECT 12.890 27.390 13.290 27.790 ;
        RECT 14.890 27.390 15.290 27.790 ;
        RECT 16.890 27.390 17.290 27.790 ;
        RECT 18.890 27.390 19.290 27.790 ;
        RECT 20.890 27.390 21.290 27.790 ;
        RECT 22.890 27.390 23.290 27.790 ;
        RECT 24.890 27.390 25.290 27.790 ;
        RECT 26.890 27.390 27.290 27.790 ;
        RECT 28.890 27.390 29.290 27.790 ;
        RECT 30.890 27.390 31.290 27.790 ;
        RECT 32.890 27.390 33.290 27.790 ;
        RECT 34.890 27.390 35.290 27.790 ;
        RECT 36.890 27.390 37.290 27.790 ;
        RECT 38.890 27.390 39.290 27.790 ;
        RECT 40.890 27.390 41.290 27.790 ;
        RECT 42.890 27.390 43.290 27.790 ;
        RECT 44.890 27.390 45.290 27.790 ;
        RECT 46.890 27.390 47.290 27.790 ;
        RECT 48.890 27.390 49.290 27.790 ;
        RECT 50.890 27.390 51.290 27.790 ;
        RECT 52.890 27.390 53.290 27.790 ;
        RECT 54.890 27.390 55.290 27.790 ;
        RECT 56.890 27.390 57.290 27.790 ;
        RECT 58.890 27.390 59.290 27.790 ;
        RECT 60.890 27.390 61.290 27.790 ;
        RECT 62.890 27.390 63.290 27.790 ;
        RECT 64.890 27.390 65.290 27.790 ;
        RECT 66.890 27.390 67.290 27.790 ;
        RECT 68.890 27.390 69.290 27.790 ;
        RECT 70.890 27.390 71.290 27.790 ;
        RECT 72.890 27.390 73.290 27.790 ;
        RECT 87.825 27.390 88.225 27.790 ;
        RECT 89.825 27.390 90.225 27.790 ;
        RECT 91.825 27.390 92.225 27.790 ;
        RECT 93.825 27.390 94.225 27.790 ;
        RECT 95.825 27.390 96.225 27.790 ;
        RECT 97.825 27.390 98.225 27.790 ;
        RECT 99.825 27.390 100.225 27.790 ;
        RECT 101.825 27.390 102.225 27.790 ;
        RECT 103.825 27.390 104.225 27.790 ;
        RECT 105.825 27.390 106.225 27.790 ;
        RECT 107.825 27.390 108.225 27.790 ;
        RECT 109.825 27.390 110.225 27.790 ;
        RECT 111.825 27.390 112.225 27.790 ;
        RECT 113.825 27.390 114.225 27.790 ;
        RECT 115.825 27.390 116.225 27.790 ;
        RECT 117.825 27.390 118.225 27.790 ;
        RECT 119.825 27.390 120.225 27.790 ;
        RECT 121.825 27.390 122.225 27.790 ;
        RECT 123.825 27.390 124.225 27.790 ;
        RECT 125.825 27.390 126.225 27.790 ;
        RECT 127.825 27.390 128.225 27.790 ;
        RECT 129.825 27.390 130.225 27.790 ;
        RECT 131.825 27.390 132.225 27.790 ;
        RECT 133.825 27.390 134.225 27.790 ;
        RECT 135.825 27.390 136.225 27.790 ;
        RECT 137.825 27.390 138.225 27.790 ;
        RECT 139.825 27.390 140.225 27.790 ;
        RECT 141.825 27.390 142.225 27.790 ;
        RECT 143.825 27.390 144.225 27.790 ;
        RECT 145.825 27.390 146.225 27.790 ;
        RECT 147.825 27.390 148.225 27.790 ;
        RECT 149.825 27.390 150.225 27.790 ;
        RECT 151.825 27.390 152.225 27.790 ;
        RECT 153.825 27.390 154.225 27.790 ;
        RECT 6.960 26.540 7.220 27.390 ;
        RECT 8.990 26.540 9.190 27.390 ;
        RECT 10.990 26.540 11.190 27.390 ;
        RECT 12.990 26.540 13.190 27.390 ;
        RECT 14.990 26.540 15.190 27.390 ;
        RECT 16.990 26.540 17.190 27.390 ;
        RECT 18.990 26.540 19.190 27.390 ;
        RECT 20.990 26.540 21.190 27.390 ;
        RECT 22.990 26.540 23.190 27.390 ;
        RECT 137.925 26.540 138.125 27.390 ;
        RECT 139.925 26.540 140.125 27.390 ;
        RECT 141.925 26.540 142.125 27.390 ;
        RECT 143.925 26.540 144.125 27.390 ;
        RECT 145.925 26.540 146.125 27.390 ;
        RECT 147.925 26.540 148.125 27.390 ;
        RECT 149.925 26.540 150.125 27.390 ;
        RECT 151.925 26.540 152.125 27.390 ;
        RECT 153.895 26.540 154.155 27.390 ;
        RECT 6.890 26.140 7.290 26.540 ;
        RECT 8.890 26.140 9.290 26.540 ;
        RECT 10.890 26.140 11.290 26.540 ;
        RECT 12.890 26.140 13.290 26.540 ;
        RECT 14.890 26.140 15.290 26.540 ;
        RECT 16.890 26.140 17.290 26.540 ;
        RECT 18.890 26.140 19.290 26.540 ;
        RECT 20.890 26.140 21.290 26.540 ;
        RECT 22.890 26.140 23.290 26.540 ;
        RECT 24.890 26.140 25.290 26.540 ;
        RECT 26.890 26.140 27.290 26.540 ;
        RECT 28.890 26.140 29.290 26.540 ;
        RECT 30.890 26.140 31.290 26.540 ;
        RECT 32.890 26.140 33.290 26.540 ;
        RECT 34.890 26.140 35.290 26.540 ;
        RECT 36.890 26.140 37.290 26.540 ;
        RECT 38.890 26.140 39.290 26.540 ;
        RECT 40.890 26.140 41.290 26.540 ;
        RECT 42.890 26.140 43.290 26.540 ;
        RECT 44.890 26.140 45.290 26.540 ;
        RECT 46.890 26.140 47.290 26.540 ;
        RECT 48.890 26.140 49.290 26.540 ;
        RECT 50.890 26.140 51.290 26.540 ;
        RECT 52.890 26.140 53.290 26.540 ;
        RECT 54.890 26.140 55.290 26.540 ;
        RECT 56.890 26.140 57.290 26.540 ;
        RECT 58.890 26.140 59.290 26.540 ;
        RECT 60.890 26.140 61.290 26.540 ;
        RECT 62.890 26.140 63.290 26.540 ;
        RECT 64.890 26.140 65.290 26.540 ;
        RECT 66.890 26.140 67.290 26.540 ;
        RECT 68.890 26.140 69.290 26.540 ;
        RECT 70.890 26.140 71.290 26.540 ;
        RECT 72.890 26.140 73.290 26.540 ;
        RECT 74.930 26.140 75.350 26.220 ;
        RECT 85.765 26.140 86.185 26.220 ;
        RECT 87.825 26.140 88.225 26.540 ;
        RECT 89.825 26.140 90.225 26.540 ;
        RECT 91.825 26.140 92.225 26.540 ;
        RECT 93.825 26.140 94.225 26.540 ;
        RECT 95.825 26.140 96.225 26.540 ;
        RECT 97.825 26.140 98.225 26.540 ;
        RECT 99.825 26.140 100.225 26.540 ;
        RECT 101.825 26.140 102.225 26.540 ;
        RECT 103.825 26.140 104.225 26.540 ;
        RECT 105.825 26.140 106.225 26.540 ;
        RECT 107.825 26.140 108.225 26.540 ;
        RECT 109.825 26.140 110.225 26.540 ;
        RECT 111.825 26.140 112.225 26.540 ;
        RECT 113.825 26.140 114.225 26.540 ;
        RECT 115.825 26.140 116.225 26.540 ;
        RECT 117.825 26.140 118.225 26.540 ;
        RECT 119.825 26.140 120.225 26.540 ;
        RECT 121.825 26.140 122.225 26.540 ;
        RECT 123.825 26.140 124.225 26.540 ;
        RECT 125.825 26.140 126.225 26.540 ;
        RECT 127.825 26.140 128.225 26.540 ;
        RECT 129.825 26.140 130.225 26.540 ;
        RECT 131.825 26.140 132.225 26.540 ;
        RECT 133.825 26.140 134.225 26.540 ;
        RECT 135.825 26.140 136.225 26.540 ;
        RECT 137.825 26.140 138.225 26.540 ;
        RECT 139.825 26.140 140.225 26.540 ;
        RECT 141.825 26.140 142.225 26.540 ;
        RECT 143.825 26.140 144.225 26.540 ;
        RECT 145.825 26.140 146.225 26.540 ;
        RECT 147.825 26.140 148.225 26.540 ;
        RECT 149.825 26.140 150.225 26.540 ;
        RECT 151.825 26.140 152.225 26.540 ;
        RECT 153.825 26.140 154.225 26.540 ;
        RECT 6.890 25.940 8.540 26.140 ;
        RECT 8.890 25.940 75.790 26.140 ;
        RECT 85.325 25.940 152.225 26.140 ;
        RECT 152.575 25.940 154.225 26.140 ;
        RECT 6.890 25.540 7.290 25.940 ;
        RECT 8.890 25.540 9.290 25.940 ;
        RECT 10.890 25.540 11.290 25.940 ;
        RECT 12.890 25.540 13.290 25.940 ;
        RECT 14.890 25.540 15.290 25.940 ;
        RECT 16.890 25.540 17.290 25.940 ;
        RECT 18.890 25.540 19.290 25.940 ;
        RECT 20.890 25.540 21.290 25.940 ;
        RECT 22.890 25.540 23.290 25.940 ;
        RECT 24.890 25.540 25.290 25.940 ;
        RECT 26.890 25.540 27.290 25.940 ;
        RECT 28.890 25.540 29.290 25.940 ;
        RECT 30.890 25.540 31.290 25.940 ;
        RECT 32.890 25.540 33.290 25.940 ;
        RECT 34.890 25.540 35.290 25.940 ;
        RECT 36.890 25.540 37.290 25.940 ;
        RECT 38.890 25.540 39.290 25.940 ;
        RECT 40.890 25.540 41.290 25.940 ;
        RECT 42.890 25.540 43.290 25.940 ;
        RECT 44.890 25.540 45.290 25.940 ;
        RECT 46.890 25.540 47.290 25.940 ;
        RECT 48.890 25.540 49.290 25.940 ;
        RECT 50.890 25.540 51.290 25.940 ;
        RECT 52.890 25.540 53.290 25.940 ;
        RECT 54.890 25.540 55.290 25.940 ;
        RECT 56.890 25.540 57.290 25.940 ;
        RECT 58.890 25.540 59.290 25.940 ;
        RECT 60.890 25.540 61.290 25.940 ;
        RECT 62.890 25.540 63.290 25.940 ;
        RECT 64.890 25.540 65.290 25.940 ;
        RECT 66.890 25.540 67.290 25.940 ;
        RECT 68.890 25.540 69.290 25.940 ;
        RECT 70.890 25.540 71.290 25.940 ;
        RECT 72.890 25.540 73.290 25.940 ;
        RECT 74.930 25.860 75.350 25.940 ;
        RECT 85.765 25.860 86.185 25.940 ;
        RECT 87.825 25.540 88.225 25.940 ;
        RECT 89.825 25.540 90.225 25.940 ;
        RECT 91.825 25.540 92.225 25.940 ;
        RECT 93.825 25.540 94.225 25.940 ;
        RECT 95.825 25.540 96.225 25.940 ;
        RECT 97.825 25.540 98.225 25.940 ;
        RECT 99.825 25.540 100.225 25.940 ;
        RECT 101.825 25.540 102.225 25.940 ;
        RECT 103.825 25.540 104.225 25.940 ;
        RECT 105.825 25.540 106.225 25.940 ;
        RECT 107.825 25.540 108.225 25.940 ;
        RECT 109.825 25.540 110.225 25.940 ;
        RECT 111.825 25.540 112.225 25.940 ;
        RECT 113.825 25.540 114.225 25.940 ;
        RECT 115.825 25.540 116.225 25.940 ;
        RECT 117.825 25.540 118.225 25.940 ;
        RECT 119.825 25.540 120.225 25.940 ;
        RECT 121.825 25.540 122.225 25.940 ;
        RECT 123.825 25.540 124.225 25.940 ;
        RECT 125.825 25.540 126.225 25.940 ;
        RECT 127.825 25.540 128.225 25.940 ;
        RECT 129.825 25.540 130.225 25.940 ;
        RECT 131.825 25.540 132.225 25.940 ;
        RECT 133.825 25.540 134.225 25.940 ;
        RECT 135.825 25.540 136.225 25.940 ;
        RECT 137.825 25.540 138.225 25.940 ;
        RECT 139.825 25.540 140.225 25.940 ;
        RECT 141.825 25.540 142.225 25.940 ;
        RECT 143.825 25.540 144.225 25.940 ;
        RECT 145.825 25.540 146.225 25.940 ;
        RECT 147.825 25.540 148.225 25.940 ;
        RECT 149.825 25.540 150.225 25.940 ;
        RECT 151.825 25.540 152.225 25.940 ;
        RECT 153.825 25.540 154.225 25.940 ;
        RECT 6.960 24.690 7.220 25.540 ;
        RECT 8.990 24.690 9.190 25.540 ;
        RECT 10.990 24.690 11.190 25.540 ;
        RECT 12.990 24.690 13.190 25.540 ;
        RECT 14.990 24.690 15.190 25.540 ;
        RECT 16.990 24.690 17.190 25.540 ;
        RECT 18.990 24.690 19.190 25.540 ;
        RECT 20.990 24.690 21.190 25.540 ;
        RECT 22.990 24.690 23.190 25.540 ;
        RECT 24.990 24.690 25.190 25.540 ;
        RECT 26.990 24.690 27.190 25.540 ;
        RECT 28.990 24.690 29.190 25.540 ;
        RECT 30.990 24.690 31.190 25.540 ;
        RECT 32.990 24.690 33.190 25.540 ;
        RECT 34.990 24.690 35.190 25.540 ;
        RECT 36.990 24.690 37.190 25.540 ;
        RECT 38.990 24.690 39.190 25.540 ;
        RECT 40.990 24.690 41.190 25.540 ;
        RECT 42.990 24.690 43.190 25.540 ;
        RECT 44.990 24.690 45.190 25.540 ;
        RECT 46.990 24.690 47.190 25.540 ;
        RECT 48.990 24.690 49.190 25.540 ;
        RECT 50.990 24.690 51.190 25.540 ;
        RECT 52.990 24.690 53.190 25.540 ;
        RECT 54.990 24.690 55.190 25.540 ;
        RECT 56.990 24.690 57.190 25.540 ;
        RECT 58.990 24.690 59.190 25.540 ;
        RECT 60.990 24.690 61.190 25.540 ;
        RECT 62.990 24.690 63.190 25.540 ;
        RECT 64.990 24.690 65.190 25.540 ;
        RECT 66.990 24.690 67.190 25.540 ;
        RECT 68.990 24.690 69.190 25.540 ;
        RECT 70.990 24.690 71.190 25.540 ;
        RECT 89.925 24.690 90.125 25.540 ;
        RECT 91.925 24.690 92.125 25.540 ;
        RECT 93.925 24.690 94.125 25.540 ;
        RECT 95.925 24.690 96.125 25.540 ;
        RECT 97.925 24.690 98.125 25.540 ;
        RECT 99.925 24.690 100.125 25.540 ;
        RECT 101.925 24.690 102.125 25.540 ;
        RECT 103.925 24.690 104.125 25.540 ;
        RECT 105.925 24.690 106.125 25.540 ;
        RECT 107.925 24.690 108.125 25.540 ;
        RECT 109.925 24.690 110.125 25.540 ;
        RECT 111.925 24.690 112.125 25.540 ;
        RECT 113.925 24.690 114.125 25.540 ;
        RECT 115.925 24.690 116.125 25.540 ;
        RECT 117.925 24.690 118.125 25.540 ;
        RECT 119.925 24.690 120.125 25.540 ;
        RECT 121.925 24.690 122.125 25.540 ;
        RECT 123.925 24.690 124.125 25.540 ;
        RECT 125.925 24.690 126.125 25.540 ;
        RECT 127.925 24.690 128.125 25.540 ;
        RECT 129.925 24.690 130.125 25.540 ;
        RECT 131.925 24.690 132.125 25.540 ;
        RECT 133.925 24.690 134.125 25.540 ;
        RECT 135.925 24.690 136.125 25.540 ;
        RECT 137.925 24.690 138.125 25.540 ;
        RECT 139.925 24.690 140.125 25.540 ;
        RECT 141.925 24.690 142.125 25.540 ;
        RECT 143.925 24.690 144.125 25.540 ;
        RECT 145.925 24.690 146.125 25.540 ;
        RECT 147.925 24.690 148.125 25.540 ;
        RECT 149.925 24.690 150.125 25.540 ;
        RECT 151.925 24.690 152.125 25.540 ;
        RECT 153.895 24.690 154.155 25.540 ;
        RECT 6.890 24.290 7.290 24.690 ;
        RECT 8.890 24.290 9.290 24.690 ;
        RECT 10.890 24.290 11.290 24.690 ;
        RECT 12.890 24.290 13.290 24.690 ;
        RECT 14.890 24.290 15.290 24.690 ;
        RECT 16.890 24.290 17.290 24.690 ;
        RECT 18.890 24.290 19.290 24.690 ;
        RECT 20.890 24.290 21.290 24.690 ;
        RECT 22.890 24.290 23.290 24.690 ;
        RECT 24.890 24.290 25.290 24.690 ;
        RECT 26.890 24.290 27.290 24.690 ;
        RECT 28.890 24.290 29.290 24.690 ;
        RECT 30.890 24.290 31.290 24.690 ;
        RECT 32.890 24.290 33.290 24.690 ;
        RECT 34.890 24.290 35.290 24.690 ;
        RECT 36.890 24.290 37.290 24.690 ;
        RECT 38.890 24.290 39.290 24.690 ;
        RECT 40.890 24.290 41.290 24.690 ;
        RECT 42.890 24.290 43.290 24.690 ;
        RECT 44.890 24.290 45.290 24.690 ;
        RECT 46.890 24.290 47.290 24.690 ;
        RECT 48.890 24.290 49.290 24.690 ;
        RECT 50.890 24.290 51.290 24.690 ;
        RECT 52.890 24.290 53.290 24.690 ;
        RECT 54.890 24.290 55.290 24.690 ;
        RECT 56.890 24.290 57.290 24.690 ;
        RECT 58.890 24.290 59.290 24.690 ;
        RECT 60.890 24.290 61.290 24.690 ;
        RECT 62.890 24.290 63.290 24.690 ;
        RECT 64.890 24.290 65.290 24.690 ;
        RECT 66.890 24.290 67.290 24.690 ;
        RECT 68.890 24.290 69.290 24.690 ;
        RECT 70.890 24.290 71.290 24.690 ;
        RECT 72.890 24.290 73.290 24.690 ;
        RECT 87.825 24.290 88.225 24.690 ;
        RECT 89.825 24.290 90.225 24.690 ;
        RECT 91.825 24.290 92.225 24.690 ;
        RECT 93.825 24.290 94.225 24.690 ;
        RECT 95.825 24.290 96.225 24.690 ;
        RECT 97.825 24.290 98.225 24.690 ;
        RECT 99.825 24.290 100.225 24.690 ;
        RECT 101.825 24.290 102.225 24.690 ;
        RECT 103.825 24.290 104.225 24.690 ;
        RECT 105.825 24.290 106.225 24.690 ;
        RECT 107.825 24.290 108.225 24.690 ;
        RECT 109.825 24.290 110.225 24.690 ;
        RECT 111.825 24.290 112.225 24.690 ;
        RECT 113.825 24.290 114.225 24.690 ;
        RECT 115.825 24.290 116.225 24.690 ;
        RECT 117.825 24.290 118.225 24.690 ;
        RECT 119.825 24.290 120.225 24.690 ;
        RECT 121.825 24.290 122.225 24.690 ;
        RECT 123.825 24.290 124.225 24.690 ;
        RECT 125.825 24.290 126.225 24.690 ;
        RECT 127.825 24.290 128.225 24.690 ;
        RECT 129.825 24.290 130.225 24.690 ;
        RECT 131.825 24.290 132.225 24.690 ;
        RECT 133.825 24.290 134.225 24.690 ;
        RECT 135.825 24.290 136.225 24.690 ;
        RECT 137.825 24.290 138.225 24.690 ;
        RECT 139.825 24.290 140.225 24.690 ;
        RECT 141.825 24.290 142.225 24.690 ;
        RECT 143.825 24.290 144.225 24.690 ;
        RECT 145.825 24.290 146.225 24.690 ;
        RECT 147.825 24.290 148.225 24.690 ;
        RECT 149.825 24.290 150.225 24.690 ;
        RECT 151.825 24.290 152.225 24.690 ;
        RECT 153.825 24.290 154.225 24.690 ;
        RECT 6.890 24.090 8.540 24.290 ;
        RECT 8.890 24.090 74.540 24.290 ;
        RECT 86.575 24.090 152.225 24.290 ;
        RECT 152.575 24.090 154.225 24.290 ;
        RECT 6.890 23.690 7.290 24.090 ;
        RECT 8.890 23.690 9.290 24.090 ;
        RECT 10.890 23.690 11.290 24.090 ;
        RECT 12.890 23.690 13.290 24.090 ;
        RECT 14.890 23.690 15.290 24.090 ;
        RECT 16.890 23.690 17.290 24.090 ;
        RECT 18.890 23.690 19.290 24.090 ;
        RECT 20.890 23.690 21.290 24.090 ;
        RECT 22.890 23.690 23.290 24.090 ;
        RECT 24.890 23.690 25.290 24.090 ;
        RECT 26.890 23.690 27.290 24.090 ;
        RECT 28.890 23.690 29.290 24.090 ;
        RECT 30.890 23.690 31.290 24.090 ;
        RECT 32.890 23.690 33.290 24.090 ;
        RECT 34.890 23.690 35.290 24.090 ;
        RECT 36.890 23.690 37.290 24.090 ;
        RECT 38.890 23.690 39.290 24.090 ;
        RECT 40.890 23.690 41.290 24.090 ;
        RECT 42.890 23.690 43.290 24.090 ;
        RECT 44.890 23.690 45.290 24.090 ;
        RECT 46.890 23.690 47.290 24.090 ;
        RECT 48.890 23.690 49.290 24.090 ;
        RECT 50.890 23.690 51.290 24.090 ;
        RECT 52.890 23.690 53.290 24.090 ;
        RECT 54.890 23.690 55.290 24.090 ;
        RECT 56.890 23.690 57.290 24.090 ;
        RECT 58.890 23.690 59.290 24.090 ;
        RECT 60.890 23.690 61.290 24.090 ;
        RECT 62.890 23.690 63.290 24.090 ;
        RECT 64.890 23.690 65.290 24.090 ;
        RECT 66.890 23.690 67.290 24.090 ;
        RECT 68.890 23.690 69.290 24.090 ;
        RECT 70.890 23.690 71.290 24.090 ;
        RECT 72.890 23.690 73.290 24.090 ;
        RECT 87.825 23.690 88.225 24.090 ;
        RECT 89.825 23.690 90.225 24.090 ;
        RECT 91.825 23.690 92.225 24.090 ;
        RECT 93.825 23.690 94.225 24.090 ;
        RECT 95.825 23.690 96.225 24.090 ;
        RECT 97.825 23.690 98.225 24.090 ;
        RECT 99.825 23.690 100.225 24.090 ;
        RECT 101.825 23.690 102.225 24.090 ;
        RECT 103.825 23.690 104.225 24.090 ;
        RECT 105.825 23.690 106.225 24.090 ;
        RECT 107.825 23.690 108.225 24.090 ;
        RECT 109.825 23.690 110.225 24.090 ;
        RECT 111.825 23.690 112.225 24.090 ;
        RECT 113.825 23.690 114.225 24.090 ;
        RECT 115.825 23.690 116.225 24.090 ;
        RECT 117.825 23.690 118.225 24.090 ;
        RECT 119.825 23.690 120.225 24.090 ;
        RECT 121.825 23.690 122.225 24.090 ;
        RECT 123.825 23.690 124.225 24.090 ;
        RECT 125.825 23.690 126.225 24.090 ;
        RECT 127.825 23.690 128.225 24.090 ;
        RECT 129.825 23.690 130.225 24.090 ;
        RECT 131.825 23.690 132.225 24.090 ;
        RECT 133.825 23.690 134.225 24.090 ;
        RECT 135.825 23.690 136.225 24.090 ;
        RECT 137.825 23.690 138.225 24.090 ;
        RECT 139.825 23.690 140.225 24.090 ;
        RECT 141.825 23.690 142.225 24.090 ;
        RECT 143.825 23.690 144.225 24.090 ;
        RECT 145.825 23.690 146.225 24.090 ;
        RECT 147.825 23.690 148.225 24.090 ;
        RECT 149.825 23.690 150.225 24.090 ;
        RECT 151.825 23.690 152.225 24.090 ;
        RECT 153.825 23.690 154.225 24.090 ;
        RECT 6.960 22.840 7.220 23.690 ;
        RECT 8.990 22.840 9.190 23.690 ;
        RECT 10.990 22.840 11.190 23.690 ;
        RECT 12.990 22.840 13.190 23.690 ;
        RECT 14.990 22.840 15.190 23.690 ;
        RECT 16.990 22.840 17.190 23.690 ;
        RECT 18.990 22.840 19.190 23.690 ;
        RECT 20.990 22.840 21.190 23.690 ;
        RECT 22.990 22.840 23.190 23.690 ;
        RECT 24.990 22.840 25.190 23.690 ;
        RECT 26.990 22.840 27.190 23.690 ;
        RECT 28.990 22.840 29.190 23.690 ;
        RECT 30.990 22.840 31.190 23.690 ;
        RECT 32.990 22.840 33.190 23.690 ;
        RECT 34.990 22.840 35.190 23.690 ;
        RECT 36.990 22.840 37.190 23.690 ;
        RECT 38.990 22.840 39.190 23.690 ;
        RECT 40.990 22.840 41.190 23.690 ;
        RECT 42.990 22.840 43.190 23.690 ;
        RECT 44.990 22.840 45.190 23.690 ;
        RECT 46.990 22.840 47.190 23.690 ;
        RECT 48.990 22.840 49.190 23.690 ;
        RECT 50.990 22.840 51.190 23.690 ;
        RECT 52.990 22.840 53.190 23.690 ;
        RECT 54.990 22.840 55.190 23.690 ;
        RECT 56.990 22.840 57.190 23.690 ;
        RECT 58.990 22.840 59.190 23.690 ;
        RECT 60.990 22.840 61.190 23.690 ;
        RECT 62.990 22.840 63.190 23.690 ;
        RECT 64.990 22.840 65.190 23.690 ;
        RECT 66.990 22.840 67.190 23.690 ;
        RECT 68.990 22.840 69.190 23.690 ;
        RECT 70.990 22.840 71.190 23.690 ;
        RECT 89.925 22.840 90.125 23.690 ;
        RECT 91.925 22.840 92.125 23.690 ;
        RECT 93.925 22.840 94.125 23.690 ;
        RECT 95.925 22.840 96.125 23.690 ;
        RECT 97.925 22.840 98.125 23.690 ;
        RECT 99.925 22.840 100.125 23.690 ;
        RECT 101.925 22.840 102.125 23.690 ;
        RECT 103.925 22.840 104.125 23.690 ;
        RECT 105.925 22.840 106.125 23.690 ;
        RECT 107.925 22.840 108.125 23.690 ;
        RECT 109.925 22.840 110.125 23.690 ;
        RECT 111.925 22.840 112.125 23.690 ;
        RECT 113.925 22.840 114.125 23.690 ;
        RECT 115.925 22.840 116.125 23.690 ;
        RECT 117.925 22.840 118.125 23.690 ;
        RECT 119.925 22.840 120.125 23.690 ;
        RECT 121.925 22.840 122.125 23.690 ;
        RECT 123.925 22.840 124.125 23.690 ;
        RECT 125.925 22.840 126.125 23.690 ;
        RECT 127.925 22.840 128.125 23.690 ;
        RECT 129.925 22.840 130.125 23.690 ;
        RECT 131.925 22.840 132.125 23.690 ;
        RECT 133.925 22.840 134.125 23.690 ;
        RECT 135.925 22.840 136.125 23.690 ;
        RECT 137.925 22.840 138.125 23.690 ;
        RECT 139.925 22.840 140.125 23.690 ;
        RECT 141.925 22.840 142.125 23.690 ;
        RECT 143.925 22.840 144.125 23.690 ;
        RECT 145.925 22.840 146.125 23.690 ;
        RECT 147.925 22.840 148.125 23.690 ;
        RECT 149.925 22.840 150.125 23.690 ;
        RECT 151.925 22.840 152.125 23.690 ;
        RECT 153.895 22.840 154.155 23.690 ;
        RECT 6.890 22.440 7.290 22.840 ;
        RECT 8.890 22.440 9.290 22.840 ;
        RECT 10.890 22.440 11.290 22.840 ;
        RECT 12.890 22.440 13.290 22.840 ;
        RECT 14.890 22.440 15.290 22.840 ;
        RECT 16.890 22.440 17.290 22.840 ;
        RECT 18.890 22.440 19.290 22.840 ;
        RECT 20.890 22.440 21.290 22.840 ;
        RECT 22.890 22.440 23.290 22.840 ;
        RECT 24.890 22.440 25.290 22.840 ;
        RECT 26.890 22.440 27.290 22.840 ;
        RECT 28.890 22.440 29.290 22.840 ;
        RECT 30.890 22.440 31.290 22.840 ;
        RECT 32.890 22.440 33.290 22.840 ;
        RECT 34.890 22.440 35.290 22.840 ;
        RECT 36.890 22.440 37.290 22.840 ;
        RECT 38.890 22.440 39.290 22.840 ;
        RECT 40.890 22.440 41.290 22.840 ;
        RECT 42.890 22.440 43.290 22.840 ;
        RECT 44.890 22.440 45.290 22.840 ;
        RECT 46.890 22.440 47.290 22.840 ;
        RECT 48.890 22.440 49.290 22.840 ;
        RECT 50.890 22.440 51.290 22.840 ;
        RECT 52.890 22.440 53.290 22.840 ;
        RECT 54.890 22.440 55.290 22.840 ;
        RECT 56.890 22.440 57.290 22.840 ;
        RECT 58.890 22.440 59.290 22.840 ;
        RECT 60.890 22.440 61.290 22.840 ;
        RECT 62.890 22.440 63.290 22.840 ;
        RECT 64.890 22.440 65.290 22.840 ;
        RECT 66.890 22.440 67.290 22.840 ;
        RECT 68.890 22.440 69.290 22.840 ;
        RECT 70.890 22.440 71.290 22.840 ;
        RECT 72.890 22.440 73.290 22.840 ;
        RECT 87.825 22.440 88.225 22.840 ;
        RECT 89.825 22.440 90.225 22.840 ;
        RECT 91.825 22.440 92.225 22.840 ;
        RECT 93.825 22.440 94.225 22.840 ;
        RECT 95.825 22.440 96.225 22.840 ;
        RECT 97.825 22.440 98.225 22.840 ;
        RECT 99.825 22.440 100.225 22.840 ;
        RECT 101.825 22.440 102.225 22.840 ;
        RECT 103.825 22.440 104.225 22.840 ;
        RECT 105.825 22.440 106.225 22.840 ;
        RECT 107.825 22.440 108.225 22.840 ;
        RECT 109.825 22.440 110.225 22.840 ;
        RECT 111.825 22.440 112.225 22.840 ;
        RECT 113.825 22.440 114.225 22.840 ;
        RECT 115.825 22.440 116.225 22.840 ;
        RECT 117.825 22.440 118.225 22.840 ;
        RECT 119.825 22.440 120.225 22.840 ;
        RECT 121.825 22.440 122.225 22.840 ;
        RECT 123.825 22.440 124.225 22.840 ;
        RECT 125.825 22.440 126.225 22.840 ;
        RECT 127.825 22.440 128.225 22.840 ;
        RECT 129.825 22.440 130.225 22.840 ;
        RECT 131.825 22.440 132.225 22.840 ;
        RECT 133.825 22.440 134.225 22.840 ;
        RECT 135.825 22.440 136.225 22.840 ;
        RECT 137.825 22.440 138.225 22.840 ;
        RECT 139.825 22.440 140.225 22.840 ;
        RECT 141.825 22.440 142.225 22.840 ;
        RECT 143.825 22.440 144.225 22.840 ;
        RECT 145.825 22.440 146.225 22.840 ;
        RECT 147.825 22.440 148.225 22.840 ;
        RECT 149.825 22.440 150.225 22.840 ;
        RECT 151.825 22.440 152.225 22.840 ;
        RECT 153.825 22.440 154.225 22.840 ;
        RECT 6.890 22.240 8.540 22.440 ;
        RECT 8.890 22.240 74.540 22.440 ;
        RECT 86.575 22.240 152.225 22.440 ;
        RECT 152.575 22.240 154.225 22.440 ;
        RECT 6.890 21.840 7.290 22.240 ;
        RECT 8.890 21.840 9.290 22.240 ;
        RECT 10.890 21.840 11.290 22.240 ;
        RECT 12.890 21.840 13.290 22.240 ;
        RECT 14.890 21.840 15.290 22.240 ;
        RECT 16.890 21.840 17.290 22.240 ;
        RECT 18.890 21.840 19.290 22.240 ;
        RECT 20.890 21.840 21.290 22.240 ;
        RECT 22.890 21.840 23.290 22.240 ;
        RECT 24.890 21.840 25.290 22.240 ;
        RECT 26.890 21.840 27.290 22.240 ;
        RECT 28.890 21.840 29.290 22.240 ;
        RECT 30.890 21.840 31.290 22.240 ;
        RECT 32.890 21.840 33.290 22.240 ;
        RECT 34.890 21.840 35.290 22.240 ;
        RECT 36.890 21.840 37.290 22.240 ;
        RECT 38.890 21.840 39.290 22.240 ;
        RECT 40.890 21.840 41.290 22.240 ;
        RECT 42.890 21.840 43.290 22.240 ;
        RECT 44.890 21.840 45.290 22.240 ;
        RECT 46.890 21.840 47.290 22.240 ;
        RECT 48.890 21.840 49.290 22.240 ;
        RECT 50.890 21.840 51.290 22.240 ;
        RECT 52.890 21.840 53.290 22.240 ;
        RECT 54.890 21.840 55.290 22.240 ;
        RECT 56.890 21.840 57.290 22.240 ;
        RECT 58.890 21.840 59.290 22.240 ;
        RECT 60.890 21.840 61.290 22.240 ;
        RECT 62.890 21.840 63.290 22.240 ;
        RECT 64.890 21.840 65.290 22.240 ;
        RECT 66.890 21.840 67.290 22.240 ;
        RECT 68.890 21.840 69.290 22.240 ;
        RECT 70.890 21.840 71.290 22.240 ;
        RECT 72.890 21.840 73.290 22.240 ;
        RECT 87.825 21.840 88.225 22.240 ;
        RECT 89.825 21.840 90.225 22.240 ;
        RECT 91.825 21.840 92.225 22.240 ;
        RECT 93.825 21.840 94.225 22.240 ;
        RECT 95.825 21.840 96.225 22.240 ;
        RECT 97.825 21.840 98.225 22.240 ;
        RECT 99.825 21.840 100.225 22.240 ;
        RECT 101.825 21.840 102.225 22.240 ;
        RECT 103.825 21.840 104.225 22.240 ;
        RECT 105.825 21.840 106.225 22.240 ;
        RECT 107.825 21.840 108.225 22.240 ;
        RECT 109.825 21.840 110.225 22.240 ;
        RECT 111.825 21.840 112.225 22.240 ;
        RECT 113.825 21.840 114.225 22.240 ;
        RECT 115.825 21.840 116.225 22.240 ;
        RECT 117.825 21.840 118.225 22.240 ;
        RECT 119.825 21.840 120.225 22.240 ;
        RECT 121.825 21.840 122.225 22.240 ;
        RECT 123.825 21.840 124.225 22.240 ;
        RECT 125.825 21.840 126.225 22.240 ;
        RECT 127.825 21.840 128.225 22.240 ;
        RECT 129.825 21.840 130.225 22.240 ;
        RECT 131.825 21.840 132.225 22.240 ;
        RECT 133.825 21.840 134.225 22.240 ;
        RECT 135.825 21.840 136.225 22.240 ;
        RECT 137.825 21.840 138.225 22.240 ;
        RECT 139.825 21.840 140.225 22.240 ;
        RECT 141.825 21.840 142.225 22.240 ;
        RECT 143.825 21.840 144.225 22.240 ;
        RECT 145.825 21.840 146.225 22.240 ;
        RECT 147.825 21.840 148.225 22.240 ;
        RECT 149.825 21.840 150.225 22.240 ;
        RECT 151.825 21.840 152.225 22.240 ;
        RECT 153.825 21.840 154.225 22.240 ;
        RECT 6.960 20.990 7.220 21.840 ;
        RECT 8.990 20.990 9.190 21.840 ;
        RECT 10.990 20.990 11.190 21.840 ;
        RECT 12.990 20.990 13.190 21.840 ;
        RECT 14.990 20.990 15.190 21.840 ;
        RECT 16.990 20.990 17.190 21.840 ;
        RECT 18.990 20.990 19.190 21.840 ;
        RECT 20.990 20.990 21.190 21.840 ;
        RECT 22.990 20.990 23.190 21.840 ;
        RECT 24.990 20.990 25.190 21.840 ;
        RECT 26.990 20.990 27.190 21.840 ;
        RECT 28.990 20.990 29.190 21.840 ;
        RECT 30.990 20.990 31.190 21.840 ;
        RECT 32.990 20.990 33.190 21.840 ;
        RECT 34.990 20.990 35.190 21.840 ;
        RECT 36.990 20.990 37.190 21.840 ;
        RECT 38.990 20.990 39.190 21.840 ;
        RECT 40.990 20.990 41.190 21.840 ;
        RECT 42.990 20.990 43.190 21.840 ;
        RECT 44.990 20.990 45.190 21.840 ;
        RECT 46.990 20.990 47.190 21.840 ;
        RECT 48.990 20.990 49.190 21.840 ;
        RECT 50.990 20.990 51.190 21.840 ;
        RECT 52.990 20.990 53.190 21.840 ;
        RECT 54.990 20.990 55.190 21.840 ;
        RECT 56.990 20.990 57.190 21.840 ;
        RECT 58.990 20.990 59.190 21.840 ;
        RECT 60.990 20.990 61.190 21.840 ;
        RECT 62.990 20.990 63.190 21.840 ;
        RECT 64.990 20.990 65.190 21.840 ;
        RECT 66.990 20.990 67.190 21.840 ;
        RECT 68.990 20.990 69.190 21.840 ;
        RECT 70.990 20.990 71.190 21.840 ;
        RECT 89.925 20.990 90.125 21.840 ;
        RECT 91.925 20.990 92.125 21.840 ;
        RECT 93.925 20.990 94.125 21.840 ;
        RECT 95.925 20.990 96.125 21.840 ;
        RECT 97.925 20.990 98.125 21.840 ;
        RECT 99.925 20.990 100.125 21.840 ;
        RECT 101.925 20.990 102.125 21.840 ;
        RECT 103.925 20.990 104.125 21.840 ;
        RECT 105.925 20.990 106.125 21.840 ;
        RECT 107.925 20.990 108.125 21.840 ;
        RECT 109.925 20.990 110.125 21.840 ;
        RECT 111.925 20.990 112.125 21.840 ;
        RECT 113.925 20.990 114.125 21.840 ;
        RECT 115.925 20.990 116.125 21.840 ;
        RECT 117.925 20.990 118.125 21.840 ;
        RECT 119.925 20.990 120.125 21.840 ;
        RECT 121.925 20.990 122.125 21.840 ;
        RECT 123.925 20.990 124.125 21.840 ;
        RECT 125.925 20.990 126.125 21.840 ;
        RECT 127.925 20.990 128.125 21.840 ;
        RECT 129.925 20.990 130.125 21.840 ;
        RECT 131.925 20.990 132.125 21.840 ;
        RECT 133.925 20.990 134.125 21.840 ;
        RECT 135.925 20.990 136.125 21.840 ;
        RECT 137.925 20.990 138.125 21.840 ;
        RECT 139.925 20.990 140.125 21.840 ;
        RECT 141.925 20.990 142.125 21.840 ;
        RECT 143.925 20.990 144.125 21.840 ;
        RECT 145.925 20.990 146.125 21.840 ;
        RECT 147.925 20.990 148.125 21.840 ;
        RECT 149.925 20.990 150.125 21.840 ;
        RECT 151.925 20.990 152.125 21.840 ;
        RECT 153.895 20.990 154.155 21.840 ;
        RECT 6.890 20.590 7.290 20.990 ;
        RECT 8.890 20.590 9.290 20.990 ;
        RECT 10.890 20.590 11.290 20.990 ;
        RECT 12.890 20.590 13.290 20.990 ;
        RECT 14.890 20.590 15.290 20.990 ;
        RECT 16.890 20.590 17.290 20.990 ;
        RECT 18.890 20.590 19.290 20.990 ;
        RECT 20.890 20.590 21.290 20.990 ;
        RECT 22.890 20.590 23.290 20.990 ;
        RECT 24.890 20.590 25.290 20.990 ;
        RECT 26.890 20.590 27.290 20.990 ;
        RECT 28.890 20.590 29.290 20.990 ;
        RECT 30.890 20.590 31.290 20.990 ;
        RECT 32.890 20.590 33.290 20.990 ;
        RECT 34.890 20.590 35.290 20.990 ;
        RECT 36.890 20.590 37.290 20.990 ;
        RECT 38.890 20.590 39.290 20.990 ;
        RECT 40.890 20.590 41.290 20.990 ;
        RECT 42.890 20.590 43.290 20.990 ;
        RECT 44.890 20.590 45.290 20.990 ;
        RECT 46.890 20.590 47.290 20.990 ;
        RECT 48.890 20.590 49.290 20.990 ;
        RECT 50.890 20.590 51.290 20.990 ;
        RECT 52.890 20.590 53.290 20.990 ;
        RECT 54.890 20.590 55.290 20.990 ;
        RECT 56.890 20.590 57.290 20.990 ;
        RECT 58.890 20.590 59.290 20.990 ;
        RECT 60.890 20.590 61.290 20.990 ;
        RECT 62.890 20.590 63.290 20.990 ;
        RECT 64.890 20.590 65.290 20.990 ;
        RECT 66.890 20.590 67.290 20.990 ;
        RECT 68.890 20.590 69.290 20.990 ;
        RECT 70.890 20.590 71.290 20.990 ;
        RECT 72.890 20.590 73.290 20.990 ;
        RECT 87.825 20.590 88.225 20.990 ;
        RECT 89.825 20.590 90.225 20.990 ;
        RECT 91.825 20.590 92.225 20.990 ;
        RECT 93.825 20.590 94.225 20.990 ;
        RECT 95.825 20.590 96.225 20.990 ;
        RECT 97.825 20.590 98.225 20.990 ;
        RECT 99.825 20.590 100.225 20.990 ;
        RECT 101.825 20.590 102.225 20.990 ;
        RECT 103.825 20.590 104.225 20.990 ;
        RECT 105.825 20.590 106.225 20.990 ;
        RECT 107.825 20.590 108.225 20.990 ;
        RECT 109.825 20.590 110.225 20.990 ;
        RECT 111.825 20.590 112.225 20.990 ;
        RECT 113.825 20.590 114.225 20.990 ;
        RECT 115.825 20.590 116.225 20.990 ;
        RECT 117.825 20.590 118.225 20.990 ;
        RECT 119.825 20.590 120.225 20.990 ;
        RECT 121.825 20.590 122.225 20.990 ;
        RECT 123.825 20.590 124.225 20.990 ;
        RECT 125.825 20.590 126.225 20.990 ;
        RECT 127.825 20.590 128.225 20.990 ;
        RECT 129.825 20.590 130.225 20.990 ;
        RECT 131.825 20.590 132.225 20.990 ;
        RECT 133.825 20.590 134.225 20.990 ;
        RECT 135.825 20.590 136.225 20.990 ;
        RECT 137.825 20.590 138.225 20.990 ;
        RECT 139.825 20.590 140.225 20.990 ;
        RECT 141.825 20.590 142.225 20.990 ;
        RECT 143.825 20.590 144.225 20.990 ;
        RECT 145.825 20.590 146.225 20.990 ;
        RECT 147.825 20.590 148.225 20.990 ;
        RECT 149.825 20.590 150.225 20.990 ;
        RECT 151.825 20.590 152.225 20.990 ;
        RECT 153.825 20.590 154.225 20.990 ;
        RECT 6.890 20.390 8.540 20.590 ;
        RECT 8.890 20.390 74.540 20.590 ;
        RECT 86.575 20.390 152.225 20.590 ;
        RECT 152.575 20.390 154.225 20.590 ;
        RECT 6.890 19.990 7.290 20.390 ;
        RECT 8.890 19.990 9.290 20.390 ;
        RECT 10.890 19.990 11.290 20.390 ;
        RECT 12.890 19.990 13.290 20.390 ;
        RECT 14.890 19.990 15.290 20.390 ;
        RECT 16.890 19.990 17.290 20.390 ;
        RECT 18.890 19.990 19.290 20.390 ;
        RECT 20.890 19.990 21.290 20.390 ;
        RECT 22.890 19.990 23.290 20.390 ;
        RECT 24.890 19.990 25.290 20.390 ;
        RECT 26.890 19.990 27.290 20.390 ;
        RECT 28.890 19.990 29.290 20.390 ;
        RECT 30.890 19.990 31.290 20.390 ;
        RECT 32.890 19.990 33.290 20.390 ;
        RECT 34.890 19.990 35.290 20.390 ;
        RECT 36.890 19.990 37.290 20.390 ;
        RECT 38.890 19.990 39.290 20.390 ;
        RECT 40.890 19.990 41.290 20.390 ;
        RECT 42.890 19.990 43.290 20.390 ;
        RECT 44.890 19.990 45.290 20.390 ;
        RECT 46.890 19.990 47.290 20.390 ;
        RECT 48.890 19.990 49.290 20.390 ;
        RECT 50.890 19.990 51.290 20.390 ;
        RECT 52.890 19.990 53.290 20.390 ;
        RECT 54.890 19.990 55.290 20.390 ;
        RECT 56.890 19.990 57.290 20.390 ;
        RECT 58.890 19.990 59.290 20.390 ;
        RECT 60.890 19.990 61.290 20.390 ;
        RECT 62.890 19.990 63.290 20.390 ;
        RECT 64.890 19.990 65.290 20.390 ;
        RECT 66.890 19.990 67.290 20.390 ;
        RECT 68.890 19.990 69.290 20.390 ;
        RECT 70.890 19.990 71.290 20.390 ;
        RECT 72.890 19.990 73.290 20.390 ;
        RECT 87.825 19.990 88.225 20.390 ;
        RECT 89.825 19.990 90.225 20.390 ;
        RECT 91.825 19.990 92.225 20.390 ;
        RECT 93.825 19.990 94.225 20.390 ;
        RECT 95.825 19.990 96.225 20.390 ;
        RECT 97.825 19.990 98.225 20.390 ;
        RECT 99.825 19.990 100.225 20.390 ;
        RECT 101.825 19.990 102.225 20.390 ;
        RECT 103.825 19.990 104.225 20.390 ;
        RECT 105.825 19.990 106.225 20.390 ;
        RECT 107.825 19.990 108.225 20.390 ;
        RECT 109.825 19.990 110.225 20.390 ;
        RECT 111.825 19.990 112.225 20.390 ;
        RECT 113.825 19.990 114.225 20.390 ;
        RECT 115.825 19.990 116.225 20.390 ;
        RECT 117.825 19.990 118.225 20.390 ;
        RECT 119.825 19.990 120.225 20.390 ;
        RECT 121.825 19.990 122.225 20.390 ;
        RECT 123.825 19.990 124.225 20.390 ;
        RECT 125.825 19.990 126.225 20.390 ;
        RECT 127.825 19.990 128.225 20.390 ;
        RECT 129.825 19.990 130.225 20.390 ;
        RECT 131.825 19.990 132.225 20.390 ;
        RECT 133.825 19.990 134.225 20.390 ;
        RECT 135.825 19.990 136.225 20.390 ;
        RECT 137.825 19.990 138.225 20.390 ;
        RECT 139.825 19.990 140.225 20.390 ;
        RECT 141.825 19.990 142.225 20.390 ;
        RECT 143.825 19.990 144.225 20.390 ;
        RECT 145.825 19.990 146.225 20.390 ;
        RECT 147.825 19.990 148.225 20.390 ;
        RECT 149.825 19.990 150.225 20.390 ;
        RECT 151.825 19.990 152.225 20.390 ;
        RECT 153.825 19.990 154.225 20.390 ;
        RECT 6.960 19.140 7.220 19.990 ;
        RECT 8.990 19.140 9.190 19.990 ;
        RECT 10.990 19.140 11.190 19.990 ;
        RECT 12.990 19.140 13.190 19.990 ;
        RECT 14.990 19.140 15.190 19.990 ;
        RECT 16.990 19.140 17.190 19.990 ;
        RECT 18.990 19.140 19.190 19.990 ;
        RECT 20.990 19.140 21.190 19.990 ;
        RECT 22.990 19.140 23.190 19.990 ;
        RECT 24.990 19.140 25.190 19.990 ;
        RECT 26.990 19.140 27.190 19.990 ;
        RECT 28.990 19.140 29.190 19.990 ;
        RECT 30.990 19.140 31.190 19.990 ;
        RECT 32.990 19.140 33.190 19.990 ;
        RECT 34.990 19.140 35.190 19.990 ;
        RECT 36.990 19.140 37.190 19.990 ;
        RECT 38.990 19.140 39.190 19.990 ;
        RECT 40.990 19.140 41.190 19.990 ;
        RECT 42.990 19.140 43.190 19.990 ;
        RECT 44.990 19.140 45.190 19.990 ;
        RECT 46.990 19.140 47.190 19.990 ;
        RECT 48.990 19.140 49.190 19.990 ;
        RECT 50.990 19.140 51.190 19.990 ;
        RECT 52.990 19.140 53.190 19.990 ;
        RECT 54.990 19.140 55.190 19.990 ;
        RECT 56.990 19.140 57.190 19.990 ;
        RECT 58.990 19.140 59.190 19.990 ;
        RECT 60.990 19.140 61.190 19.990 ;
        RECT 62.990 19.140 63.190 19.990 ;
        RECT 64.990 19.140 65.190 19.990 ;
        RECT 66.990 19.140 67.190 19.990 ;
        RECT 68.990 19.140 69.190 19.990 ;
        RECT 70.990 19.140 71.190 19.990 ;
        RECT 89.925 19.140 90.125 19.990 ;
        RECT 91.925 19.140 92.125 19.990 ;
        RECT 93.925 19.140 94.125 19.990 ;
        RECT 95.925 19.140 96.125 19.990 ;
        RECT 97.925 19.140 98.125 19.990 ;
        RECT 99.925 19.140 100.125 19.990 ;
        RECT 101.925 19.140 102.125 19.990 ;
        RECT 103.925 19.140 104.125 19.990 ;
        RECT 105.925 19.140 106.125 19.990 ;
        RECT 107.925 19.140 108.125 19.990 ;
        RECT 109.925 19.140 110.125 19.990 ;
        RECT 111.925 19.140 112.125 19.990 ;
        RECT 113.925 19.140 114.125 19.990 ;
        RECT 115.925 19.140 116.125 19.990 ;
        RECT 117.925 19.140 118.125 19.990 ;
        RECT 119.925 19.140 120.125 19.990 ;
        RECT 121.925 19.140 122.125 19.990 ;
        RECT 123.925 19.140 124.125 19.990 ;
        RECT 125.925 19.140 126.125 19.990 ;
        RECT 127.925 19.140 128.125 19.990 ;
        RECT 129.925 19.140 130.125 19.990 ;
        RECT 131.925 19.140 132.125 19.990 ;
        RECT 133.925 19.140 134.125 19.990 ;
        RECT 135.925 19.140 136.125 19.990 ;
        RECT 137.925 19.140 138.125 19.990 ;
        RECT 139.925 19.140 140.125 19.990 ;
        RECT 141.925 19.140 142.125 19.990 ;
        RECT 143.925 19.140 144.125 19.990 ;
        RECT 145.925 19.140 146.125 19.990 ;
        RECT 147.925 19.140 148.125 19.990 ;
        RECT 149.925 19.140 150.125 19.990 ;
        RECT 151.925 19.140 152.125 19.990 ;
        RECT 153.895 19.140 154.155 19.990 ;
        RECT 6.890 18.740 7.290 19.140 ;
        RECT 8.890 18.740 9.290 19.140 ;
        RECT 10.890 18.740 11.290 19.140 ;
        RECT 12.890 18.740 13.290 19.140 ;
        RECT 14.890 18.740 15.290 19.140 ;
        RECT 16.890 18.740 17.290 19.140 ;
        RECT 18.890 18.740 19.290 19.140 ;
        RECT 20.890 18.740 21.290 19.140 ;
        RECT 22.890 18.740 23.290 19.140 ;
        RECT 24.890 18.740 25.290 19.140 ;
        RECT 26.890 18.740 27.290 19.140 ;
        RECT 28.890 18.740 29.290 19.140 ;
        RECT 30.890 18.740 31.290 19.140 ;
        RECT 32.890 18.740 33.290 19.140 ;
        RECT 34.890 18.740 35.290 19.140 ;
        RECT 36.890 18.740 37.290 19.140 ;
        RECT 38.890 18.740 39.290 19.140 ;
        RECT 40.890 18.740 41.290 19.140 ;
        RECT 42.890 18.740 43.290 19.140 ;
        RECT 44.890 18.740 45.290 19.140 ;
        RECT 46.890 18.740 47.290 19.140 ;
        RECT 48.890 18.740 49.290 19.140 ;
        RECT 50.890 18.740 51.290 19.140 ;
        RECT 52.890 18.740 53.290 19.140 ;
        RECT 54.890 18.740 55.290 19.140 ;
        RECT 56.890 18.740 57.290 19.140 ;
        RECT 58.890 18.740 59.290 19.140 ;
        RECT 60.890 18.740 61.290 19.140 ;
        RECT 62.890 18.740 63.290 19.140 ;
        RECT 64.890 18.740 65.290 19.140 ;
        RECT 66.890 18.740 67.290 19.140 ;
        RECT 68.890 18.740 69.290 19.140 ;
        RECT 70.890 18.740 71.290 19.140 ;
        RECT 72.890 18.740 73.290 19.140 ;
        RECT 87.825 18.740 88.225 19.140 ;
        RECT 89.825 18.740 90.225 19.140 ;
        RECT 91.825 18.740 92.225 19.140 ;
        RECT 93.825 18.740 94.225 19.140 ;
        RECT 95.825 18.740 96.225 19.140 ;
        RECT 97.825 18.740 98.225 19.140 ;
        RECT 99.825 18.740 100.225 19.140 ;
        RECT 101.825 18.740 102.225 19.140 ;
        RECT 103.825 18.740 104.225 19.140 ;
        RECT 105.825 18.740 106.225 19.140 ;
        RECT 107.825 18.740 108.225 19.140 ;
        RECT 109.825 18.740 110.225 19.140 ;
        RECT 111.825 18.740 112.225 19.140 ;
        RECT 113.825 18.740 114.225 19.140 ;
        RECT 115.825 18.740 116.225 19.140 ;
        RECT 117.825 18.740 118.225 19.140 ;
        RECT 119.825 18.740 120.225 19.140 ;
        RECT 121.825 18.740 122.225 19.140 ;
        RECT 123.825 18.740 124.225 19.140 ;
        RECT 125.825 18.740 126.225 19.140 ;
        RECT 127.825 18.740 128.225 19.140 ;
        RECT 129.825 18.740 130.225 19.140 ;
        RECT 131.825 18.740 132.225 19.140 ;
        RECT 133.825 18.740 134.225 19.140 ;
        RECT 135.825 18.740 136.225 19.140 ;
        RECT 137.825 18.740 138.225 19.140 ;
        RECT 139.825 18.740 140.225 19.140 ;
        RECT 141.825 18.740 142.225 19.140 ;
        RECT 143.825 18.740 144.225 19.140 ;
        RECT 145.825 18.740 146.225 19.140 ;
        RECT 147.825 18.740 148.225 19.140 ;
        RECT 149.825 18.740 150.225 19.140 ;
        RECT 151.825 18.740 152.225 19.140 ;
        RECT 153.825 18.740 154.225 19.140 ;
        RECT 6.890 18.540 8.540 18.740 ;
        RECT 8.890 18.540 74.540 18.740 ;
        RECT 86.575 18.540 152.225 18.740 ;
        RECT 152.575 18.540 154.225 18.740 ;
        RECT 6.890 18.140 7.290 18.540 ;
        RECT 8.890 18.140 9.290 18.540 ;
        RECT 10.890 18.140 11.290 18.540 ;
        RECT 12.890 18.140 13.290 18.540 ;
        RECT 14.890 18.140 15.290 18.540 ;
        RECT 16.890 18.140 17.290 18.540 ;
        RECT 18.890 18.140 19.290 18.540 ;
        RECT 20.890 18.140 21.290 18.540 ;
        RECT 22.890 18.140 23.290 18.540 ;
        RECT 24.890 18.140 25.290 18.540 ;
        RECT 26.890 18.140 27.290 18.540 ;
        RECT 28.890 18.140 29.290 18.540 ;
        RECT 30.890 18.140 31.290 18.540 ;
        RECT 32.890 18.140 33.290 18.540 ;
        RECT 34.890 18.140 35.290 18.540 ;
        RECT 36.890 18.140 37.290 18.540 ;
        RECT 38.890 18.140 39.290 18.540 ;
        RECT 40.890 18.140 41.290 18.540 ;
        RECT 42.890 18.140 43.290 18.540 ;
        RECT 44.890 18.140 45.290 18.540 ;
        RECT 46.890 18.140 47.290 18.540 ;
        RECT 48.890 18.140 49.290 18.540 ;
        RECT 50.890 18.140 51.290 18.540 ;
        RECT 52.890 18.140 53.290 18.540 ;
        RECT 54.890 18.140 55.290 18.540 ;
        RECT 56.890 18.140 57.290 18.540 ;
        RECT 58.890 18.140 59.290 18.540 ;
        RECT 60.890 18.140 61.290 18.540 ;
        RECT 62.890 18.140 63.290 18.540 ;
        RECT 64.890 18.140 65.290 18.540 ;
        RECT 66.890 18.140 67.290 18.540 ;
        RECT 68.890 18.140 69.290 18.540 ;
        RECT 70.890 18.140 71.290 18.540 ;
        RECT 72.890 18.140 73.290 18.540 ;
        RECT 87.825 18.140 88.225 18.540 ;
        RECT 89.825 18.140 90.225 18.540 ;
        RECT 91.825 18.140 92.225 18.540 ;
        RECT 93.825 18.140 94.225 18.540 ;
        RECT 95.825 18.140 96.225 18.540 ;
        RECT 97.825 18.140 98.225 18.540 ;
        RECT 99.825 18.140 100.225 18.540 ;
        RECT 101.825 18.140 102.225 18.540 ;
        RECT 103.825 18.140 104.225 18.540 ;
        RECT 105.825 18.140 106.225 18.540 ;
        RECT 107.825 18.140 108.225 18.540 ;
        RECT 109.825 18.140 110.225 18.540 ;
        RECT 111.825 18.140 112.225 18.540 ;
        RECT 113.825 18.140 114.225 18.540 ;
        RECT 115.825 18.140 116.225 18.540 ;
        RECT 117.825 18.140 118.225 18.540 ;
        RECT 119.825 18.140 120.225 18.540 ;
        RECT 121.825 18.140 122.225 18.540 ;
        RECT 123.825 18.140 124.225 18.540 ;
        RECT 125.825 18.140 126.225 18.540 ;
        RECT 127.825 18.140 128.225 18.540 ;
        RECT 129.825 18.140 130.225 18.540 ;
        RECT 131.825 18.140 132.225 18.540 ;
        RECT 133.825 18.140 134.225 18.540 ;
        RECT 135.825 18.140 136.225 18.540 ;
        RECT 137.825 18.140 138.225 18.540 ;
        RECT 139.825 18.140 140.225 18.540 ;
        RECT 141.825 18.140 142.225 18.540 ;
        RECT 143.825 18.140 144.225 18.540 ;
        RECT 145.825 18.140 146.225 18.540 ;
        RECT 147.825 18.140 148.225 18.540 ;
        RECT 149.825 18.140 150.225 18.540 ;
        RECT 151.825 18.140 152.225 18.540 ;
        RECT 153.825 18.140 154.225 18.540 ;
        RECT 6.960 17.290 7.220 18.140 ;
        RECT 8.990 17.290 9.190 18.140 ;
        RECT 10.990 17.290 11.190 18.140 ;
        RECT 12.990 17.290 13.190 18.140 ;
        RECT 14.990 17.290 15.190 18.140 ;
        RECT 16.990 17.290 17.190 18.140 ;
        RECT 18.990 17.290 19.190 18.140 ;
        RECT 20.990 17.290 21.190 18.140 ;
        RECT 22.990 17.290 23.190 18.140 ;
        RECT 24.990 17.290 25.190 18.140 ;
        RECT 26.990 17.290 27.190 18.140 ;
        RECT 28.990 17.290 29.190 18.140 ;
        RECT 30.990 17.290 31.190 18.140 ;
        RECT 32.990 17.290 33.190 18.140 ;
        RECT 34.990 17.290 35.190 18.140 ;
        RECT 36.990 17.290 37.190 18.140 ;
        RECT 38.990 17.290 39.190 18.140 ;
        RECT 40.990 17.290 41.190 18.140 ;
        RECT 42.990 17.290 43.190 18.140 ;
        RECT 44.990 17.290 45.190 18.140 ;
        RECT 46.990 17.290 47.190 18.140 ;
        RECT 48.990 17.290 49.190 18.140 ;
        RECT 50.990 17.290 51.190 18.140 ;
        RECT 52.990 17.290 53.190 18.140 ;
        RECT 54.990 17.290 55.190 18.140 ;
        RECT 56.990 17.290 57.190 18.140 ;
        RECT 58.990 17.290 59.190 18.140 ;
        RECT 60.990 17.290 61.190 18.140 ;
        RECT 62.990 17.290 63.190 18.140 ;
        RECT 64.990 17.290 65.190 18.140 ;
        RECT 66.990 17.290 67.190 18.140 ;
        RECT 68.990 17.290 69.190 18.140 ;
        RECT 70.990 17.290 71.190 18.140 ;
        RECT 89.925 17.290 90.125 18.140 ;
        RECT 91.925 17.290 92.125 18.140 ;
        RECT 93.925 17.290 94.125 18.140 ;
        RECT 95.925 17.290 96.125 18.140 ;
        RECT 97.925 17.290 98.125 18.140 ;
        RECT 99.925 17.290 100.125 18.140 ;
        RECT 101.925 17.290 102.125 18.140 ;
        RECT 103.925 17.290 104.125 18.140 ;
        RECT 105.925 17.290 106.125 18.140 ;
        RECT 107.925 17.290 108.125 18.140 ;
        RECT 109.925 17.290 110.125 18.140 ;
        RECT 111.925 17.290 112.125 18.140 ;
        RECT 113.925 17.290 114.125 18.140 ;
        RECT 115.925 17.290 116.125 18.140 ;
        RECT 117.925 17.290 118.125 18.140 ;
        RECT 119.925 17.290 120.125 18.140 ;
        RECT 121.925 17.290 122.125 18.140 ;
        RECT 123.925 17.290 124.125 18.140 ;
        RECT 125.925 17.290 126.125 18.140 ;
        RECT 127.925 17.290 128.125 18.140 ;
        RECT 129.925 17.290 130.125 18.140 ;
        RECT 131.925 17.290 132.125 18.140 ;
        RECT 133.925 17.290 134.125 18.140 ;
        RECT 135.925 17.290 136.125 18.140 ;
        RECT 137.925 17.290 138.125 18.140 ;
        RECT 139.925 17.290 140.125 18.140 ;
        RECT 141.925 17.290 142.125 18.140 ;
        RECT 143.925 17.290 144.125 18.140 ;
        RECT 145.925 17.290 146.125 18.140 ;
        RECT 147.925 17.290 148.125 18.140 ;
        RECT 149.925 17.290 150.125 18.140 ;
        RECT 151.925 17.290 152.125 18.140 ;
        RECT 153.895 17.290 154.155 18.140 ;
        RECT 6.890 16.890 7.290 17.290 ;
        RECT 8.890 16.890 9.290 17.290 ;
        RECT 10.890 16.890 11.290 17.290 ;
        RECT 12.890 16.890 13.290 17.290 ;
        RECT 14.890 16.890 15.290 17.290 ;
        RECT 16.890 16.890 17.290 17.290 ;
        RECT 18.890 16.890 19.290 17.290 ;
        RECT 20.890 16.890 21.290 17.290 ;
        RECT 22.890 16.890 23.290 17.290 ;
        RECT 24.890 16.890 25.290 17.290 ;
        RECT 26.890 16.890 27.290 17.290 ;
        RECT 28.890 16.890 29.290 17.290 ;
        RECT 30.890 16.890 31.290 17.290 ;
        RECT 32.890 16.890 33.290 17.290 ;
        RECT 34.890 16.890 35.290 17.290 ;
        RECT 36.890 16.890 37.290 17.290 ;
        RECT 38.890 16.890 39.290 17.290 ;
        RECT 40.890 16.890 41.290 17.290 ;
        RECT 42.890 16.890 43.290 17.290 ;
        RECT 44.890 16.890 45.290 17.290 ;
        RECT 46.890 16.890 47.290 17.290 ;
        RECT 48.890 16.890 49.290 17.290 ;
        RECT 50.890 16.890 51.290 17.290 ;
        RECT 52.890 16.890 53.290 17.290 ;
        RECT 54.890 16.890 55.290 17.290 ;
        RECT 56.890 16.890 57.290 17.290 ;
        RECT 58.890 16.890 59.290 17.290 ;
        RECT 60.890 16.890 61.290 17.290 ;
        RECT 62.890 16.890 63.290 17.290 ;
        RECT 64.890 16.890 65.290 17.290 ;
        RECT 66.890 16.890 67.290 17.290 ;
        RECT 68.890 16.890 69.290 17.290 ;
        RECT 70.890 16.890 71.290 17.290 ;
        RECT 72.890 16.890 73.290 17.290 ;
        RECT 87.825 16.890 88.225 17.290 ;
        RECT 89.825 16.890 90.225 17.290 ;
        RECT 91.825 16.890 92.225 17.290 ;
        RECT 93.825 16.890 94.225 17.290 ;
        RECT 95.825 16.890 96.225 17.290 ;
        RECT 97.825 16.890 98.225 17.290 ;
        RECT 99.825 16.890 100.225 17.290 ;
        RECT 101.825 16.890 102.225 17.290 ;
        RECT 103.825 16.890 104.225 17.290 ;
        RECT 105.825 16.890 106.225 17.290 ;
        RECT 107.825 16.890 108.225 17.290 ;
        RECT 109.825 16.890 110.225 17.290 ;
        RECT 111.825 16.890 112.225 17.290 ;
        RECT 113.825 16.890 114.225 17.290 ;
        RECT 115.825 16.890 116.225 17.290 ;
        RECT 117.825 16.890 118.225 17.290 ;
        RECT 119.825 16.890 120.225 17.290 ;
        RECT 121.825 16.890 122.225 17.290 ;
        RECT 123.825 16.890 124.225 17.290 ;
        RECT 125.825 16.890 126.225 17.290 ;
        RECT 127.825 16.890 128.225 17.290 ;
        RECT 129.825 16.890 130.225 17.290 ;
        RECT 131.825 16.890 132.225 17.290 ;
        RECT 133.825 16.890 134.225 17.290 ;
        RECT 135.825 16.890 136.225 17.290 ;
        RECT 137.825 16.890 138.225 17.290 ;
        RECT 139.825 16.890 140.225 17.290 ;
        RECT 141.825 16.890 142.225 17.290 ;
        RECT 143.825 16.890 144.225 17.290 ;
        RECT 145.825 16.890 146.225 17.290 ;
        RECT 147.825 16.890 148.225 17.290 ;
        RECT 149.825 16.890 150.225 17.290 ;
        RECT 151.825 16.890 152.225 17.290 ;
        RECT 153.825 16.890 154.225 17.290 ;
        RECT 6.890 16.690 8.540 16.890 ;
        RECT 8.890 16.690 74.540 16.890 ;
        RECT 86.575 16.690 152.225 16.890 ;
        RECT 152.575 16.690 154.225 16.890 ;
        RECT 6.890 16.290 7.290 16.690 ;
        RECT 8.890 16.290 9.290 16.690 ;
        RECT 10.890 16.290 11.290 16.690 ;
        RECT 12.890 16.290 13.290 16.690 ;
        RECT 14.890 16.290 15.290 16.690 ;
        RECT 16.890 16.290 17.290 16.690 ;
        RECT 18.890 16.290 19.290 16.690 ;
        RECT 20.890 16.290 21.290 16.690 ;
        RECT 22.890 16.290 23.290 16.690 ;
        RECT 24.890 16.290 25.290 16.690 ;
        RECT 26.890 16.290 27.290 16.690 ;
        RECT 28.890 16.290 29.290 16.690 ;
        RECT 30.890 16.290 31.290 16.690 ;
        RECT 32.890 16.290 33.290 16.690 ;
        RECT 34.890 16.290 35.290 16.690 ;
        RECT 36.890 16.290 37.290 16.690 ;
        RECT 38.890 16.290 39.290 16.690 ;
        RECT 40.890 16.290 41.290 16.690 ;
        RECT 42.890 16.290 43.290 16.690 ;
        RECT 44.890 16.290 45.290 16.690 ;
        RECT 46.890 16.290 47.290 16.690 ;
        RECT 48.890 16.290 49.290 16.690 ;
        RECT 50.890 16.290 51.290 16.690 ;
        RECT 52.890 16.290 53.290 16.690 ;
        RECT 54.890 16.290 55.290 16.690 ;
        RECT 56.890 16.290 57.290 16.690 ;
        RECT 58.890 16.290 59.290 16.690 ;
        RECT 60.890 16.290 61.290 16.690 ;
        RECT 62.890 16.290 63.290 16.690 ;
        RECT 64.890 16.290 65.290 16.690 ;
        RECT 66.890 16.290 67.290 16.690 ;
        RECT 68.890 16.290 69.290 16.690 ;
        RECT 70.890 16.290 71.290 16.690 ;
        RECT 72.890 16.290 73.290 16.690 ;
        RECT 87.825 16.290 88.225 16.690 ;
        RECT 89.825 16.290 90.225 16.690 ;
        RECT 91.825 16.290 92.225 16.690 ;
        RECT 93.825 16.290 94.225 16.690 ;
        RECT 95.825 16.290 96.225 16.690 ;
        RECT 97.825 16.290 98.225 16.690 ;
        RECT 99.825 16.290 100.225 16.690 ;
        RECT 101.825 16.290 102.225 16.690 ;
        RECT 103.825 16.290 104.225 16.690 ;
        RECT 105.825 16.290 106.225 16.690 ;
        RECT 107.825 16.290 108.225 16.690 ;
        RECT 109.825 16.290 110.225 16.690 ;
        RECT 111.825 16.290 112.225 16.690 ;
        RECT 113.825 16.290 114.225 16.690 ;
        RECT 115.825 16.290 116.225 16.690 ;
        RECT 117.825 16.290 118.225 16.690 ;
        RECT 119.825 16.290 120.225 16.690 ;
        RECT 121.825 16.290 122.225 16.690 ;
        RECT 123.825 16.290 124.225 16.690 ;
        RECT 125.825 16.290 126.225 16.690 ;
        RECT 127.825 16.290 128.225 16.690 ;
        RECT 129.825 16.290 130.225 16.690 ;
        RECT 131.825 16.290 132.225 16.690 ;
        RECT 133.825 16.290 134.225 16.690 ;
        RECT 135.825 16.290 136.225 16.690 ;
        RECT 137.825 16.290 138.225 16.690 ;
        RECT 139.825 16.290 140.225 16.690 ;
        RECT 141.825 16.290 142.225 16.690 ;
        RECT 143.825 16.290 144.225 16.690 ;
        RECT 145.825 16.290 146.225 16.690 ;
        RECT 147.825 16.290 148.225 16.690 ;
        RECT 149.825 16.290 150.225 16.690 ;
        RECT 151.825 16.290 152.225 16.690 ;
        RECT 153.825 16.290 154.225 16.690 ;
        RECT 6.960 15.440 7.220 16.290 ;
        RECT 8.990 15.440 9.190 16.290 ;
        RECT 10.990 15.440 11.190 16.290 ;
        RECT 12.990 15.440 13.190 16.290 ;
        RECT 14.990 15.440 15.190 16.290 ;
        RECT 16.990 15.440 17.190 16.290 ;
        RECT 18.990 15.440 19.190 16.290 ;
        RECT 20.990 15.440 21.190 16.290 ;
        RECT 22.990 15.440 23.190 16.290 ;
        RECT 24.990 15.440 25.190 16.290 ;
        RECT 26.990 15.440 27.190 16.290 ;
        RECT 28.990 15.440 29.190 16.290 ;
        RECT 30.990 15.440 31.190 16.290 ;
        RECT 32.990 15.440 33.190 16.290 ;
        RECT 34.990 15.440 35.190 16.290 ;
        RECT 36.990 15.440 37.190 16.290 ;
        RECT 38.990 15.440 39.190 16.290 ;
        RECT 40.990 15.440 41.190 16.290 ;
        RECT 42.990 15.440 43.190 16.290 ;
        RECT 44.990 15.440 45.190 16.290 ;
        RECT 46.990 15.440 47.190 16.290 ;
        RECT 48.990 15.440 49.190 16.290 ;
        RECT 50.990 15.440 51.190 16.290 ;
        RECT 52.990 15.440 53.190 16.290 ;
        RECT 54.990 15.440 55.190 16.290 ;
        RECT 56.990 15.440 57.190 16.290 ;
        RECT 58.990 15.440 59.190 16.290 ;
        RECT 60.990 15.440 61.190 16.290 ;
        RECT 62.990 15.440 63.190 16.290 ;
        RECT 64.990 15.440 65.190 16.290 ;
        RECT 66.990 15.440 67.190 16.290 ;
        RECT 68.990 15.440 69.190 16.290 ;
        RECT 70.990 15.440 71.190 16.290 ;
        RECT 89.925 15.440 90.125 16.290 ;
        RECT 91.925 15.440 92.125 16.290 ;
        RECT 93.925 15.440 94.125 16.290 ;
        RECT 95.925 15.440 96.125 16.290 ;
        RECT 97.925 15.440 98.125 16.290 ;
        RECT 99.925 15.440 100.125 16.290 ;
        RECT 101.925 15.440 102.125 16.290 ;
        RECT 103.925 15.440 104.125 16.290 ;
        RECT 105.925 15.440 106.125 16.290 ;
        RECT 107.925 15.440 108.125 16.290 ;
        RECT 109.925 15.440 110.125 16.290 ;
        RECT 111.925 15.440 112.125 16.290 ;
        RECT 113.925 15.440 114.125 16.290 ;
        RECT 115.925 15.440 116.125 16.290 ;
        RECT 117.925 15.440 118.125 16.290 ;
        RECT 119.925 15.440 120.125 16.290 ;
        RECT 121.925 15.440 122.125 16.290 ;
        RECT 123.925 15.440 124.125 16.290 ;
        RECT 125.925 15.440 126.125 16.290 ;
        RECT 127.925 15.440 128.125 16.290 ;
        RECT 129.925 15.440 130.125 16.290 ;
        RECT 131.925 15.440 132.125 16.290 ;
        RECT 133.925 15.440 134.125 16.290 ;
        RECT 135.925 15.440 136.125 16.290 ;
        RECT 137.925 15.440 138.125 16.290 ;
        RECT 139.925 15.440 140.125 16.290 ;
        RECT 141.925 15.440 142.125 16.290 ;
        RECT 143.925 15.440 144.125 16.290 ;
        RECT 145.925 15.440 146.125 16.290 ;
        RECT 147.925 15.440 148.125 16.290 ;
        RECT 149.925 15.440 150.125 16.290 ;
        RECT 151.925 15.440 152.125 16.290 ;
        RECT 153.895 15.440 154.155 16.290 ;
        RECT 6.890 15.040 7.290 15.440 ;
        RECT 8.890 15.040 9.290 15.440 ;
        RECT 10.890 15.040 11.290 15.440 ;
        RECT 12.890 15.040 13.290 15.440 ;
        RECT 14.890 15.040 15.290 15.440 ;
        RECT 16.890 15.040 17.290 15.440 ;
        RECT 18.890 15.040 19.290 15.440 ;
        RECT 20.890 15.040 21.290 15.440 ;
        RECT 22.890 15.040 23.290 15.440 ;
        RECT 24.890 15.040 25.290 15.440 ;
        RECT 26.890 15.040 27.290 15.440 ;
        RECT 28.890 15.040 29.290 15.440 ;
        RECT 30.890 15.040 31.290 15.440 ;
        RECT 32.890 15.040 33.290 15.440 ;
        RECT 34.890 15.040 35.290 15.440 ;
        RECT 36.890 15.040 37.290 15.440 ;
        RECT 38.890 15.040 39.290 15.440 ;
        RECT 40.890 15.040 41.290 15.440 ;
        RECT 42.890 15.040 43.290 15.440 ;
        RECT 44.890 15.040 45.290 15.440 ;
        RECT 46.890 15.040 47.290 15.440 ;
        RECT 48.890 15.040 49.290 15.440 ;
        RECT 50.890 15.040 51.290 15.440 ;
        RECT 52.890 15.040 53.290 15.440 ;
        RECT 54.890 15.040 55.290 15.440 ;
        RECT 56.890 15.040 57.290 15.440 ;
        RECT 58.890 15.040 59.290 15.440 ;
        RECT 60.890 15.040 61.290 15.440 ;
        RECT 62.890 15.040 63.290 15.440 ;
        RECT 64.890 15.040 65.290 15.440 ;
        RECT 66.890 15.040 67.290 15.440 ;
        RECT 68.890 15.040 69.290 15.440 ;
        RECT 70.890 15.040 71.290 15.440 ;
        RECT 72.890 15.040 73.290 15.440 ;
        RECT 87.825 15.040 88.225 15.440 ;
        RECT 89.825 15.040 90.225 15.440 ;
        RECT 91.825 15.040 92.225 15.440 ;
        RECT 93.825 15.040 94.225 15.440 ;
        RECT 95.825 15.040 96.225 15.440 ;
        RECT 97.825 15.040 98.225 15.440 ;
        RECT 99.825 15.040 100.225 15.440 ;
        RECT 101.825 15.040 102.225 15.440 ;
        RECT 103.825 15.040 104.225 15.440 ;
        RECT 105.825 15.040 106.225 15.440 ;
        RECT 107.825 15.040 108.225 15.440 ;
        RECT 109.825 15.040 110.225 15.440 ;
        RECT 111.825 15.040 112.225 15.440 ;
        RECT 113.825 15.040 114.225 15.440 ;
        RECT 115.825 15.040 116.225 15.440 ;
        RECT 117.825 15.040 118.225 15.440 ;
        RECT 119.825 15.040 120.225 15.440 ;
        RECT 121.825 15.040 122.225 15.440 ;
        RECT 123.825 15.040 124.225 15.440 ;
        RECT 125.825 15.040 126.225 15.440 ;
        RECT 127.825 15.040 128.225 15.440 ;
        RECT 129.825 15.040 130.225 15.440 ;
        RECT 131.825 15.040 132.225 15.440 ;
        RECT 133.825 15.040 134.225 15.440 ;
        RECT 135.825 15.040 136.225 15.440 ;
        RECT 137.825 15.040 138.225 15.440 ;
        RECT 139.825 15.040 140.225 15.440 ;
        RECT 141.825 15.040 142.225 15.440 ;
        RECT 143.825 15.040 144.225 15.440 ;
        RECT 145.825 15.040 146.225 15.440 ;
        RECT 147.825 15.040 148.225 15.440 ;
        RECT 149.825 15.040 150.225 15.440 ;
        RECT 151.825 15.040 152.225 15.440 ;
        RECT 153.825 15.040 154.225 15.440 ;
        RECT 6.890 14.840 8.540 15.040 ;
        RECT 8.890 14.840 74.540 15.040 ;
        RECT 86.575 14.840 152.225 15.040 ;
        RECT 152.575 14.840 154.225 15.040 ;
        RECT 6.890 14.440 7.290 14.840 ;
        RECT 8.890 14.440 9.290 14.840 ;
        RECT 10.890 14.440 11.290 14.840 ;
        RECT 12.890 14.440 13.290 14.840 ;
        RECT 14.890 14.440 15.290 14.840 ;
        RECT 16.890 14.440 17.290 14.840 ;
        RECT 18.890 14.440 19.290 14.840 ;
        RECT 20.890 14.440 21.290 14.840 ;
        RECT 22.890 14.440 23.290 14.840 ;
        RECT 24.890 14.440 25.290 14.840 ;
        RECT 26.890 14.440 27.290 14.840 ;
        RECT 28.890 14.440 29.290 14.840 ;
        RECT 30.890 14.440 31.290 14.840 ;
        RECT 32.890 14.440 33.290 14.840 ;
        RECT 34.890 14.440 35.290 14.840 ;
        RECT 36.890 14.440 37.290 14.840 ;
        RECT 38.890 14.440 39.290 14.840 ;
        RECT 40.890 14.440 41.290 14.840 ;
        RECT 42.890 14.440 43.290 14.840 ;
        RECT 44.890 14.440 45.290 14.840 ;
        RECT 46.890 14.440 47.290 14.840 ;
        RECT 48.890 14.440 49.290 14.840 ;
        RECT 50.890 14.440 51.290 14.840 ;
        RECT 52.890 14.440 53.290 14.840 ;
        RECT 54.890 14.440 55.290 14.840 ;
        RECT 56.890 14.440 57.290 14.840 ;
        RECT 58.890 14.440 59.290 14.840 ;
        RECT 60.890 14.440 61.290 14.840 ;
        RECT 62.890 14.440 63.290 14.840 ;
        RECT 64.890 14.440 65.290 14.840 ;
        RECT 66.890 14.440 67.290 14.840 ;
        RECT 68.890 14.440 69.290 14.840 ;
        RECT 70.890 14.440 71.290 14.840 ;
        RECT 72.890 14.440 73.290 14.840 ;
        RECT 87.825 14.440 88.225 14.840 ;
        RECT 89.825 14.440 90.225 14.840 ;
        RECT 91.825 14.440 92.225 14.840 ;
        RECT 93.825 14.440 94.225 14.840 ;
        RECT 95.825 14.440 96.225 14.840 ;
        RECT 97.825 14.440 98.225 14.840 ;
        RECT 99.825 14.440 100.225 14.840 ;
        RECT 101.825 14.440 102.225 14.840 ;
        RECT 103.825 14.440 104.225 14.840 ;
        RECT 105.825 14.440 106.225 14.840 ;
        RECT 107.825 14.440 108.225 14.840 ;
        RECT 109.825 14.440 110.225 14.840 ;
        RECT 111.825 14.440 112.225 14.840 ;
        RECT 113.825 14.440 114.225 14.840 ;
        RECT 115.825 14.440 116.225 14.840 ;
        RECT 117.825 14.440 118.225 14.840 ;
        RECT 119.825 14.440 120.225 14.840 ;
        RECT 121.825 14.440 122.225 14.840 ;
        RECT 123.825 14.440 124.225 14.840 ;
        RECT 125.825 14.440 126.225 14.840 ;
        RECT 127.825 14.440 128.225 14.840 ;
        RECT 129.825 14.440 130.225 14.840 ;
        RECT 131.825 14.440 132.225 14.840 ;
        RECT 133.825 14.440 134.225 14.840 ;
        RECT 135.825 14.440 136.225 14.840 ;
        RECT 137.825 14.440 138.225 14.840 ;
        RECT 139.825 14.440 140.225 14.840 ;
        RECT 141.825 14.440 142.225 14.840 ;
        RECT 143.825 14.440 144.225 14.840 ;
        RECT 145.825 14.440 146.225 14.840 ;
        RECT 147.825 14.440 148.225 14.840 ;
        RECT 149.825 14.440 150.225 14.840 ;
        RECT 151.825 14.440 152.225 14.840 ;
        RECT 153.825 14.440 154.225 14.840 ;
        RECT 6.960 13.590 7.220 14.440 ;
        RECT 8.990 13.590 9.190 14.440 ;
        RECT 10.990 13.590 11.190 14.440 ;
        RECT 12.990 13.590 13.190 14.440 ;
        RECT 14.990 13.590 15.190 14.440 ;
        RECT 16.990 13.590 17.190 14.440 ;
        RECT 18.990 13.590 19.190 14.440 ;
        RECT 20.990 13.590 21.190 14.440 ;
        RECT 22.990 13.590 23.190 14.440 ;
        RECT 24.990 13.590 25.190 14.440 ;
        RECT 26.990 13.590 27.190 14.440 ;
        RECT 28.990 13.590 29.190 14.440 ;
        RECT 30.990 13.590 31.190 14.440 ;
        RECT 32.990 13.590 33.190 14.440 ;
        RECT 34.990 13.590 35.190 14.440 ;
        RECT 36.990 13.590 37.190 14.440 ;
        RECT 38.990 13.590 39.190 14.440 ;
        RECT 40.990 13.590 41.190 14.440 ;
        RECT 42.990 13.590 43.190 14.440 ;
        RECT 44.990 13.590 45.190 14.440 ;
        RECT 46.990 13.590 47.190 14.440 ;
        RECT 48.990 13.590 49.190 14.440 ;
        RECT 50.990 13.590 51.190 14.440 ;
        RECT 52.990 13.590 53.190 14.440 ;
        RECT 54.990 13.590 55.190 14.440 ;
        RECT 56.990 13.590 57.190 14.440 ;
        RECT 58.990 13.590 59.190 14.440 ;
        RECT 60.990 13.590 61.190 14.440 ;
        RECT 62.990 13.590 63.190 14.440 ;
        RECT 64.990 13.590 65.190 14.440 ;
        RECT 66.990 13.590 67.190 14.440 ;
        RECT 68.990 13.590 69.190 14.440 ;
        RECT 70.990 13.590 71.190 14.440 ;
        RECT 89.925 13.590 90.125 14.440 ;
        RECT 91.925 13.590 92.125 14.440 ;
        RECT 93.925 13.590 94.125 14.440 ;
        RECT 95.925 13.590 96.125 14.440 ;
        RECT 97.925 13.590 98.125 14.440 ;
        RECT 99.925 13.590 100.125 14.440 ;
        RECT 101.925 13.590 102.125 14.440 ;
        RECT 103.925 13.590 104.125 14.440 ;
        RECT 105.925 13.590 106.125 14.440 ;
        RECT 107.925 13.590 108.125 14.440 ;
        RECT 109.925 13.590 110.125 14.440 ;
        RECT 111.925 13.590 112.125 14.440 ;
        RECT 113.925 13.590 114.125 14.440 ;
        RECT 115.925 13.590 116.125 14.440 ;
        RECT 117.925 13.590 118.125 14.440 ;
        RECT 119.925 13.590 120.125 14.440 ;
        RECT 121.925 13.590 122.125 14.440 ;
        RECT 123.925 13.590 124.125 14.440 ;
        RECT 125.925 13.590 126.125 14.440 ;
        RECT 127.925 13.590 128.125 14.440 ;
        RECT 129.925 13.590 130.125 14.440 ;
        RECT 131.925 13.590 132.125 14.440 ;
        RECT 133.925 13.590 134.125 14.440 ;
        RECT 135.925 13.590 136.125 14.440 ;
        RECT 137.925 13.590 138.125 14.440 ;
        RECT 139.925 13.590 140.125 14.440 ;
        RECT 141.925 13.590 142.125 14.440 ;
        RECT 143.925 13.590 144.125 14.440 ;
        RECT 145.925 13.590 146.125 14.440 ;
        RECT 147.925 13.590 148.125 14.440 ;
        RECT 149.925 13.590 150.125 14.440 ;
        RECT 151.925 13.590 152.125 14.440 ;
        RECT 153.895 13.590 154.155 14.440 ;
        RECT 6.890 13.190 7.290 13.590 ;
        RECT 8.890 13.190 9.290 13.590 ;
        RECT 10.890 13.190 11.290 13.590 ;
        RECT 12.890 13.190 13.290 13.590 ;
        RECT 14.890 13.190 15.290 13.590 ;
        RECT 16.890 13.190 17.290 13.590 ;
        RECT 18.890 13.190 19.290 13.590 ;
        RECT 20.890 13.190 21.290 13.590 ;
        RECT 22.890 13.190 23.290 13.590 ;
        RECT 24.890 13.190 25.290 13.590 ;
        RECT 26.890 13.190 27.290 13.590 ;
        RECT 28.890 13.190 29.290 13.590 ;
        RECT 30.890 13.190 31.290 13.590 ;
        RECT 32.890 13.190 33.290 13.590 ;
        RECT 34.890 13.190 35.290 13.590 ;
        RECT 36.890 13.190 37.290 13.590 ;
        RECT 38.890 13.190 39.290 13.590 ;
        RECT 40.890 13.190 41.290 13.590 ;
        RECT 42.890 13.190 43.290 13.590 ;
        RECT 44.890 13.190 45.290 13.590 ;
        RECT 46.890 13.190 47.290 13.590 ;
        RECT 48.890 13.190 49.290 13.590 ;
        RECT 50.890 13.190 51.290 13.590 ;
        RECT 52.890 13.190 53.290 13.590 ;
        RECT 54.890 13.190 55.290 13.590 ;
        RECT 56.890 13.190 57.290 13.590 ;
        RECT 58.890 13.190 59.290 13.590 ;
        RECT 60.890 13.190 61.290 13.590 ;
        RECT 62.890 13.190 63.290 13.590 ;
        RECT 64.890 13.190 65.290 13.590 ;
        RECT 66.890 13.190 67.290 13.590 ;
        RECT 68.890 13.190 69.290 13.590 ;
        RECT 70.890 13.190 71.290 13.590 ;
        RECT 72.890 13.190 73.290 13.590 ;
        RECT 87.825 13.190 88.225 13.590 ;
        RECT 89.825 13.190 90.225 13.590 ;
        RECT 91.825 13.190 92.225 13.590 ;
        RECT 93.825 13.190 94.225 13.590 ;
        RECT 95.825 13.190 96.225 13.590 ;
        RECT 97.825 13.190 98.225 13.590 ;
        RECT 99.825 13.190 100.225 13.590 ;
        RECT 101.825 13.190 102.225 13.590 ;
        RECT 103.825 13.190 104.225 13.590 ;
        RECT 105.825 13.190 106.225 13.590 ;
        RECT 107.825 13.190 108.225 13.590 ;
        RECT 109.825 13.190 110.225 13.590 ;
        RECT 111.825 13.190 112.225 13.590 ;
        RECT 113.825 13.190 114.225 13.590 ;
        RECT 115.825 13.190 116.225 13.590 ;
        RECT 117.825 13.190 118.225 13.590 ;
        RECT 119.825 13.190 120.225 13.590 ;
        RECT 121.825 13.190 122.225 13.590 ;
        RECT 123.825 13.190 124.225 13.590 ;
        RECT 125.825 13.190 126.225 13.590 ;
        RECT 127.825 13.190 128.225 13.590 ;
        RECT 129.825 13.190 130.225 13.590 ;
        RECT 131.825 13.190 132.225 13.590 ;
        RECT 133.825 13.190 134.225 13.590 ;
        RECT 135.825 13.190 136.225 13.590 ;
        RECT 137.825 13.190 138.225 13.590 ;
        RECT 139.825 13.190 140.225 13.590 ;
        RECT 141.825 13.190 142.225 13.590 ;
        RECT 143.825 13.190 144.225 13.590 ;
        RECT 145.825 13.190 146.225 13.590 ;
        RECT 147.825 13.190 148.225 13.590 ;
        RECT 149.825 13.190 150.225 13.590 ;
        RECT 151.825 13.190 152.225 13.590 ;
        RECT 153.825 13.190 154.225 13.590 ;
        RECT 6.890 12.990 8.540 13.190 ;
        RECT 8.890 12.990 74.540 13.190 ;
        RECT 86.575 12.990 152.225 13.190 ;
        RECT 152.575 12.990 154.225 13.190 ;
        RECT 6.890 12.590 7.290 12.990 ;
        RECT 8.890 12.590 9.290 12.990 ;
        RECT 10.890 12.590 11.290 12.990 ;
        RECT 12.890 12.590 13.290 12.990 ;
        RECT 14.890 12.590 15.290 12.990 ;
        RECT 16.890 12.590 17.290 12.990 ;
        RECT 18.890 12.590 19.290 12.990 ;
        RECT 20.890 12.590 21.290 12.990 ;
        RECT 22.890 12.590 23.290 12.990 ;
        RECT 24.890 12.590 25.290 12.990 ;
        RECT 26.890 12.590 27.290 12.990 ;
        RECT 28.890 12.590 29.290 12.990 ;
        RECT 30.890 12.590 31.290 12.990 ;
        RECT 32.890 12.590 33.290 12.990 ;
        RECT 34.890 12.590 35.290 12.990 ;
        RECT 36.890 12.590 37.290 12.990 ;
        RECT 38.890 12.590 39.290 12.990 ;
        RECT 40.890 12.590 41.290 12.990 ;
        RECT 42.890 12.590 43.290 12.990 ;
        RECT 44.890 12.590 45.290 12.990 ;
        RECT 46.890 12.590 47.290 12.990 ;
        RECT 48.890 12.590 49.290 12.990 ;
        RECT 50.890 12.590 51.290 12.990 ;
        RECT 52.890 12.590 53.290 12.990 ;
        RECT 54.890 12.590 55.290 12.990 ;
        RECT 56.890 12.590 57.290 12.990 ;
        RECT 58.890 12.590 59.290 12.990 ;
        RECT 60.890 12.590 61.290 12.990 ;
        RECT 62.890 12.590 63.290 12.990 ;
        RECT 64.890 12.590 65.290 12.990 ;
        RECT 66.890 12.590 67.290 12.990 ;
        RECT 68.890 12.590 69.290 12.990 ;
        RECT 70.890 12.590 71.290 12.990 ;
        RECT 72.890 12.590 73.290 12.990 ;
        RECT 87.825 12.590 88.225 12.990 ;
        RECT 89.825 12.590 90.225 12.990 ;
        RECT 91.825 12.590 92.225 12.990 ;
        RECT 93.825 12.590 94.225 12.990 ;
        RECT 95.825 12.590 96.225 12.990 ;
        RECT 97.825 12.590 98.225 12.990 ;
        RECT 99.825 12.590 100.225 12.990 ;
        RECT 101.825 12.590 102.225 12.990 ;
        RECT 103.825 12.590 104.225 12.990 ;
        RECT 105.825 12.590 106.225 12.990 ;
        RECT 107.825 12.590 108.225 12.990 ;
        RECT 109.825 12.590 110.225 12.990 ;
        RECT 111.825 12.590 112.225 12.990 ;
        RECT 113.825 12.590 114.225 12.990 ;
        RECT 115.825 12.590 116.225 12.990 ;
        RECT 117.825 12.590 118.225 12.990 ;
        RECT 119.825 12.590 120.225 12.990 ;
        RECT 121.825 12.590 122.225 12.990 ;
        RECT 123.825 12.590 124.225 12.990 ;
        RECT 125.825 12.590 126.225 12.990 ;
        RECT 127.825 12.590 128.225 12.990 ;
        RECT 129.825 12.590 130.225 12.990 ;
        RECT 131.825 12.590 132.225 12.990 ;
        RECT 133.825 12.590 134.225 12.990 ;
        RECT 135.825 12.590 136.225 12.990 ;
        RECT 137.825 12.590 138.225 12.990 ;
        RECT 139.825 12.590 140.225 12.990 ;
        RECT 141.825 12.590 142.225 12.990 ;
        RECT 143.825 12.590 144.225 12.990 ;
        RECT 145.825 12.590 146.225 12.990 ;
        RECT 147.825 12.590 148.225 12.990 ;
        RECT 149.825 12.590 150.225 12.990 ;
        RECT 151.825 12.590 152.225 12.990 ;
        RECT 153.825 12.590 154.225 12.990 ;
        RECT 6.960 11.740 7.220 12.590 ;
        RECT 8.990 11.740 9.190 12.590 ;
        RECT 10.990 11.740 11.190 12.590 ;
        RECT 12.990 11.740 13.190 12.590 ;
        RECT 14.990 11.740 15.190 12.590 ;
        RECT 16.990 11.740 17.190 12.590 ;
        RECT 18.990 11.740 19.190 12.590 ;
        RECT 20.990 11.740 21.190 12.590 ;
        RECT 22.990 11.740 23.190 12.590 ;
        RECT 24.990 11.740 25.190 12.590 ;
        RECT 26.990 11.740 27.190 12.590 ;
        RECT 28.990 11.740 29.190 12.590 ;
        RECT 30.990 11.740 31.190 12.590 ;
        RECT 32.990 11.740 33.190 12.590 ;
        RECT 34.990 11.740 35.190 12.590 ;
        RECT 36.990 11.740 37.190 12.590 ;
        RECT 38.990 11.740 39.190 12.590 ;
        RECT 40.990 11.740 41.190 12.590 ;
        RECT 42.990 11.740 43.190 12.590 ;
        RECT 44.990 11.740 45.190 12.590 ;
        RECT 46.990 11.740 47.190 12.590 ;
        RECT 48.990 11.740 49.190 12.590 ;
        RECT 50.990 11.740 51.190 12.590 ;
        RECT 52.990 11.740 53.190 12.590 ;
        RECT 54.990 11.740 55.190 12.590 ;
        RECT 56.990 11.740 57.190 12.590 ;
        RECT 58.990 11.740 59.190 12.590 ;
        RECT 60.990 11.740 61.190 12.590 ;
        RECT 62.990 11.740 63.190 12.590 ;
        RECT 64.990 11.740 65.190 12.590 ;
        RECT 66.990 11.740 67.190 12.590 ;
        RECT 68.990 11.740 69.190 12.590 ;
        RECT 70.990 11.740 71.190 12.590 ;
        RECT 89.925 11.740 90.125 12.590 ;
        RECT 91.925 11.740 92.125 12.590 ;
        RECT 93.925 11.740 94.125 12.590 ;
        RECT 95.925 11.740 96.125 12.590 ;
        RECT 97.925 11.740 98.125 12.590 ;
        RECT 99.925 11.740 100.125 12.590 ;
        RECT 101.925 11.740 102.125 12.590 ;
        RECT 103.925 11.740 104.125 12.590 ;
        RECT 105.925 11.740 106.125 12.590 ;
        RECT 107.925 11.740 108.125 12.590 ;
        RECT 109.925 11.740 110.125 12.590 ;
        RECT 111.925 11.740 112.125 12.590 ;
        RECT 113.925 11.740 114.125 12.590 ;
        RECT 115.925 11.740 116.125 12.590 ;
        RECT 117.925 11.740 118.125 12.590 ;
        RECT 119.925 11.740 120.125 12.590 ;
        RECT 121.925 11.740 122.125 12.590 ;
        RECT 123.925 11.740 124.125 12.590 ;
        RECT 125.925 11.740 126.125 12.590 ;
        RECT 127.925 11.740 128.125 12.590 ;
        RECT 129.925 11.740 130.125 12.590 ;
        RECT 131.925 11.740 132.125 12.590 ;
        RECT 133.925 11.740 134.125 12.590 ;
        RECT 135.925 11.740 136.125 12.590 ;
        RECT 137.925 11.740 138.125 12.590 ;
        RECT 139.925 11.740 140.125 12.590 ;
        RECT 141.925 11.740 142.125 12.590 ;
        RECT 143.925 11.740 144.125 12.590 ;
        RECT 145.925 11.740 146.125 12.590 ;
        RECT 147.925 11.740 148.125 12.590 ;
        RECT 149.925 11.740 150.125 12.590 ;
        RECT 151.925 11.740 152.125 12.590 ;
        RECT 153.895 11.740 154.155 12.590 ;
        RECT 6.890 11.340 7.290 11.740 ;
        RECT 8.890 11.340 9.290 11.740 ;
        RECT 10.890 11.340 11.290 11.740 ;
        RECT 12.890 11.340 13.290 11.740 ;
        RECT 14.890 11.340 15.290 11.740 ;
        RECT 16.890 11.340 17.290 11.740 ;
        RECT 18.890 11.340 19.290 11.740 ;
        RECT 20.890 11.340 21.290 11.740 ;
        RECT 22.890 11.340 23.290 11.740 ;
        RECT 24.890 11.340 25.290 11.740 ;
        RECT 26.890 11.340 27.290 11.740 ;
        RECT 28.890 11.340 29.290 11.740 ;
        RECT 30.890 11.340 31.290 11.740 ;
        RECT 32.890 11.340 33.290 11.740 ;
        RECT 34.890 11.340 35.290 11.740 ;
        RECT 36.890 11.340 37.290 11.740 ;
        RECT 38.890 11.340 39.290 11.740 ;
        RECT 40.890 11.340 41.290 11.740 ;
        RECT 42.890 11.340 43.290 11.740 ;
        RECT 44.890 11.340 45.290 11.740 ;
        RECT 46.890 11.340 47.290 11.740 ;
        RECT 48.890 11.340 49.290 11.740 ;
        RECT 50.890 11.340 51.290 11.740 ;
        RECT 52.890 11.340 53.290 11.740 ;
        RECT 54.890 11.340 55.290 11.740 ;
        RECT 56.890 11.340 57.290 11.740 ;
        RECT 58.890 11.340 59.290 11.740 ;
        RECT 60.890 11.340 61.290 11.740 ;
        RECT 62.890 11.340 63.290 11.740 ;
        RECT 64.890 11.340 65.290 11.740 ;
        RECT 66.890 11.340 67.290 11.740 ;
        RECT 68.890 11.340 69.290 11.740 ;
        RECT 70.890 11.340 71.290 11.740 ;
        RECT 72.890 11.340 73.290 11.740 ;
        RECT 87.825 11.340 88.225 11.740 ;
        RECT 89.825 11.340 90.225 11.740 ;
        RECT 91.825 11.340 92.225 11.740 ;
        RECT 93.825 11.340 94.225 11.740 ;
        RECT 95.825 11.340 96.225 11.740 ;
        RECT 97.825 11.340 98.225 11.740 ;
        RECT 99.825 11.340 100.225 11.740 ;
        RECT 101.825 11.340 102.225 11.740 ;
        RECT 103.825 11.340 104.225 11.740 ;
        RECT 105.825 11.340 106.225 11.740 ;
        RECT 107.825 11.340 108.225 11.740 ;
        RECT 109.825 11.340 110.225 11.740 ;
        RECT 111.825 11.340 112.225 11.740 ;
        RECT 113.825 11.340 114.225 11.740 ;
        RECT 115.825 11.340 116.225 11.740 ;
        RECT 117.825 11.340 118.225 11.740 ;
        RECT 119.825 11.340 120.225 11.740 ;
        RECT 121.825 11.340 122.225 11.740 ;
        RECT 123.825 11.340 124.225 11.740 ;
        RECT 125.825 11.340 126.225 11.740 ;
        RECT 127.825 11.340 128.225 11.740 ;
        RECT 129.825 11.340 130.225 11.740 ;
        RECT 131.825 11.340 132.225 11.740 ;
        RECT 133.825 11.340 134.225 11.740 ;
        RECT 135.825 11.340 136.225 11.740 ;
        RECT 137.825 11.340 138.225 11.740 ;
        RECT 139.825 11.340 140.225 11.740 ;
        RECT 141.825 11.340 142.225 11.740 ;
        RECT 143.825 11.340 144.225 11.740 ;
        RECT 145.825 11.340 146.225 11.740 ;
        RECT 147.825 11.340 148.225 11.740 ;
        RECT 149.825 11.340 150.225 11.740 ;
        RECT 151.825 11.340 152.225 11.740 ;
        RECT 153.825 11.340 154.225 11.740 ;
        RECT 6.890 11.140 8.540 11.340 ;
        RECT 8.890 11.140 74.540 11.340 ;
        RECT 86.575 11.140 152.225 11.340 ;
        RECT 152.575 11.140 154.225 11.340 ;
        RECT 6.890 10.740 7.290 11.140 ;
        RECT 8.890 10.740 9.290 11.140 ;
        RECT 10.890 10.740 11.290 11.140 ;
        RECT 12.890 10.740 13.290 11.140 ;
        RECT 14.890 10.740 15.290 11.140 ;
        RECT 16.890 10.740 17.290 11.140 ;
        RECT 18.890 10.740 19.290 11.140 ;
        RECT 20.890 10.740 21.290 11.140 ;
        RECT 22.890 10.740 23.290 11.140 ;
        RECT 24.890 10.740 25.290 11.140 ;
        RECT 26.890 10.740 27.290 11.140 ;
        RECT 28.890 10.740 29.290 11.140 ;
        RECT 30.890 10.740 31.290 11.140 ;
        RECT 32.890 10.740 33.290 11.140 ;
        RECT 34.890 10.740 35.290 11.140 ;
        RECT 36.890 10.740 37.290 11.140 ;
        RECT 38.890 10.740 39.290 11.140 ;
        RECT 40.890 10.740 41.290 11.140 ;
        RECT 42.890 10.740 43.290 11.140 ;
        RECT 44.890 10.740 45.290 11.140 ;
        RECT 46.890 10.740 47.290 11.140 ;
        RECT 48.890 10.740 49.290 11.140 ;
        RECT 50.890 10.740 51.290 11.140 ;
        RECT 52.890 10.740 53.290 11.140 ;
        RECT 54.890 10.740 55.290 11.140 ;
        RECT 56.890 10.740 57.290 11.140 ;
        RECT 58.890 10.740 59.290 11.140 ;
        RECT 60.890 10.740 61.290 11.140 ;
        RECT 62.890 10.740 63.290 11.140 ;
        RECT 64.890 10.740 65.290 11.140 ;
        RECT 66.890 10.740 67.290 11.140 ;
        RECT 68.890 10.740 69.290 11.140 ;
        RECT 70.890 10.740 71.290 11.140 ;
        RECT 72.890 10.740 73.290 11.140 ;
        RECT 87.825 10.740 88.225 11.140 ;
        RECT 89.825 10.740 90.225 11.140 ;
        RECT 91.825 10.740 92.225 11.140 ;
        RECT 93.825 10.740 94.225 11.140 ;
        RECT 95.825 10.740 96.225 11.140 ;
        RECT 97.825 10.740 98.225 11.140 ;
        RECT 99.825 10.740 100.225 11.140 ;
        RECT 101.825 10.740 102.225 11.140 ;
        RECT 103.825 10.740 104.225 11.140 ;
        RECT 105.825 10.740 106.225 11.140 ;
        RECT 107.825 10.740 108.225 11.140 ;
        RECT 109.825 10.740 110.225 11.140 ;
        RECT 111.825 10.740 112.225 11.140 ;
        RECT 113.825 10.740 114.225 11.140 ;
        RECT 115.825 10.740 116.225 11.140 ;
        RECT 117.825 10.740 118.225 11.140 ;
        RECT 119.825 10.740 120.225 11.140 ;
        RECT 121.825 10.740 122.225 11.140 ;
        RECT 123.825 10.740 124.225 11.140 ;
        RECT 125.825 10.740 126.225 11.140 ;
        RECT 127.825 10.740 128.225 11.140 ;
        RECT 129.825 10.740 130.225 11.140 ;
        RECT 131.825 10.740 132.225 11.140 ;
        RECT 133.825 10.740 134.225 11.140 ;
        RECT 135.825 10.740 136.225 11.140 ;
        RECT 137.825 10.740 138.225 11.140 ;
        RECT 139.825 10.740 140.225 11.140 ;
        RECT 141.825 10.740 142.225 11.140 ;
        RECT 143.825 10.740 144.225 11.140 ;
        RECT 145.825 10.740 146.225 11.140 ;
        RECT 147.825 10.740 148.225 11.140 ;
        RECT 149.825 10.740 150.225 11.140 ;
        RECT 151.825 10.740 152.225 11.140 ;
        RECT 153.825 10.740 154.225 11.140 ;
        RECT 6.960 9.890 7.220 10.740 ;
        RECT 8.990 9.890 9.190 10.740 ;
        RECT 10.990 9.890 11.190 10.740 ;
        RECT 12.990 9.890 13.190 10.740 ;
        RECT 14.990 9.890 15.190 10.740 ;
        RECT 16.990 9.890 17.190 10.740 ;
        RECT 18.990 9.890 19.190 10.740 ;
        RECT 20.990 9.890 21.190 10.740 ;
        RECT 22.990 9.890 23.190 10.740 ;
        RECT 24.990 9.890 25.190 10.740 ;
        RECT 26.990 9.890 27.190 10.740 ;
        RECT 28.990 9.890 29.190 10.740 ;
        RECT 30.990 9.890 31.190 10.740 ;
        RECT 32.990 9.890 33.190 10.740 ;
        RECT 34.990 9.890 35.190 10.740 ;
        RECT 36.990 9.890 37.190 10.740 ;
        RECT 38.990 9.890 39.190 10.740 ;
        RECT 40.990 9.890 41.190 10.740 ;
        RECT 42.990 9.890 43.190 10.740 ;
        RECT 44.990 9.890 45.190 10.740 ;
        RECT 46.990 9.890 47.190 10.740 ;
        RECT 48.990 9.890 49.190 10.740 ;
        RECT 50.990 9.890 51.190 10.740 ;
        RECT 52.990 9.890 53.190 10.740 ;
        RECT 54.990 9.890 55.190 10.740 ;
        RECT 56.990 9.890 57.190 10.740 ;
        RECT 58.990 9.890 59.190 10.740 ;
        RECT 60.990 9.890 61.190 10.740 ;
        RECT 62.990 9.890 63.190 10.740 ;
        RECT 64.990 9.890 65.190 10.740 ;
        RECT 66.990 9.890 67.190 10.740 ;
        RECT 68.990 9.890 69.190 10.740 ;
        RECT 70.990 9.890 71.190 10.740 ;
        RECT 89.925 9.890 90.125 10.740 ;
        RECT 91.925 9.890 92.125 10.740 ;
        RECT 93.925 9.890 94.125 10.740 ;
        RECT 95.925 9.890 96.125 10.740 ;
        RECT 97.925 9.890 98.125 10.740 ;
        RECT 99.925 9.890 100.125 10.740 ;
        RECT 101.925 9.890 102.125 10.740 ;
        RECT 103.925 9.890 104.125 10.740 ;
        RECT 105.925 9.890 106.125 10.740 ;
        RECT 107.925 9.890 108.125 10.740 ;
        RECT 109.925 9.890 110.125 10.740 ;
        RECT 111.925 9.890 112.125 10.740 ;
        RECT 113.925 9.890 114.125 10.740 ;
        RECT 115.925 9.890 116.125 10.740 ;
        RECT 117.925 9.890 118.125 10.740 ;
        RECT 119.925 9.890 120.125 10.740 ;
        RECT 121.925 9.890 122.125 10.740 ;
        RECT 123.925 9.890 124.125 10.740 ;
        RECT 125.925 9.890 126.125 10.740 ;
        RECT 127.925 9.890 128.125 10.740 ;
        RECT 129.925 9.890 130.125 10.740 ;
        RECT 131.925 9.890 132.125 10.740 ;
        RECT 133.925 9.890 134.125 10.740 ;
        RECT 135.925 9.890 136.125 10.740 ;
        RECT 137.925 9.890 138.125 10.740 ;
        RECT 139.925 9.890 140.125 10.740 ;
        RECT 141.925 9.890 142.125 10.740 ;
        RECT 143.925 9.890 144.125 10.740 ;
        RECT 145.925 9.890 146.125 10.740 ;
        RECT 147.925 9.890 148.125 10.740 ;
        RECT 149.925 9.890 150.125 10.740 ;
        RECT 151.925 9.890 152.125 10.740 ;
        RECT 153.895 9.890 154.155 10.740 ;
        RECT 6.890 9.490 7.290 9.890 ;
        RECT 8.890 9.490 9.290 9.890 ;
        RECT 10.890 9.490 11.290 9.890 ;
        RECT 12.890 9.490 13.290 9.890 ;
        RECT 14.890 9.490 15.290 9.890 ;
        RECT 16.890 9.490 17.290 9.890 ;
        RECT 18.890 9.490 19.290 9.890 ;
        RECT 20.890 9.490 21.290 9.890 ;
        RECT 22.890 9.490 23.290 9.890 ;
        RECT 24.890 9.490 25.290 9.890 ;
        RECT 26.890 9.490 27.290 9.890 ;
        RECT 28.890 9.490 29.290 9.890 ;
        RECT 30.890 9.490 31.290 9.890 ;
        RECT 32.890 9.490 33.290 9.890 ;
        RECT 34.890 9.490 35.290 9.890 ;
        RECT 36.890 9.490 37.290 9.890 ;
        RECT 38.890 9.490 39.290 9.890 ;
        RECT 40.890 9.490 41.290 9.890 ;
        RECT 42.890 9.490 43.290 9.890 ;
        RECT 44.890 9.490 45.290 9.890 ;
        RECT 46.890 9.490 47.290 9.890 ;
        RECT 48.890 9.490 49.290 9.890 ;
        RECT 50.890 9.490 51.290 9.890 ;
        RECT 52.890 9.490 53.290 9.890 ;
        RECT 54.890 9.490 55.290 9.890 ;
        RECT 56.890 9.490 57.290 9.890 ;
        RECT 58.890 9.490 59.290 9.890 ;
        RECT 60.890 9.490 61.290 9.890 ;
        RECT 62.890 9.490 63.290 9.890 ;
        RECT 64.890 9.490 65.290 9.890 ;
        RECT 66.890 9.490 67.290 9.890 ;
        RECT 68.890 9.490 69.290 9.890 ;
        RECT 70.890 9.490 71.290 9.890 ;
        RECT 72.890 9.490 73.290 9.890 ;
        RECT 87.825 9.490 88.225 9.890 ;
        RECT 89.825 9.490 90.225 9.890 ;
        RECT 91.825 9.490 92.225 9.890 ;
        RECT 93.825 9.490 94.225 9.890 ;
        RECT 95.825 9.490 96.225 9.890 ;
        RECT 97.825 9.490 98.225 9.890 ;
        RECT 99.825 9.490 100.225 9.890 ;
        RECT 101.825 9.490 102.225 9.890 ;
        RECT 103.825 9.490 104.225 9.890 ;
        RECT 105.825 9.490 106.225 9.890 ;
        RECT 107.825 9.490 108.225 9.890 ;
        RECT 109.825 9.490 110.225 9.890 ;
        RECT 111.825 9.490 112.225 9.890 ;
        RECT 113.825 9.490 114.225 9.890 ;
        RECT 115.825 9.490 116.225 9.890 ;
        RECT 117.825 9.490 118.225 9.890 ;
        RECT 119.825 9.490 120.225 9.890 ;
        RECT 121.825 9.490 122.225 9.890 ;
        RECT 123.825 9.490 124.225 9.890 ;
        RECT 125.825 9.490 126.225 9.890 ;
        RECT 127.825 9.490 128.225 9.890 ;
        RECT 129.825 9.490 130.225 9.890 ;
        RECT 131.825 9.490 132.225 9.890 ;
        RECT 133.825 9.490 134.225 9.890 ;
        RECT 135.825 9.490 136.225 9.890 ;
        RECT 137.825 9.490 138.225 9.890 ;
        RECT 139.825 9.490 140.225 9.890 ;
        RECT 141.825 9.490 142.225 9.890 ;
        RECT 143.825 9.490 144.225 9.890 ;
        RECT 145.825 9.490 146.225 9.890 ;
        RECT 147.825 9.490 148.225 9.890 ;
        RECT 149.825 9.490 150.225 9.890 ;
        RECT 151.825 9.490 152.225 9.890 ;
        RECT 153.825 9.490 154.225 9.890 ;
        RECT 6.890 9.290 8.540 9.490 ;
        RECT 8.890 9.290 74.540 9.490 ;
        RECT 86.575 9.290 152.225 9.490 ;
        RECT 152.575 9.290 154.225 9.490 ;
        RECT 6.890 8.890 7.290 9.290 ;
        RECT 8.890 8.890 9.290 9.290 ;
        RECT 10.890 8.890 11.290 9.290 ;
        RECT 12.890 8.890 13.290 9.290 ;
        RECT 14.890 8.890 15.290 9.290 ;
        RECT 16.890 8.890 17.290 9.290 ;
        RECT 18.890 8.890 19.290 9.290 ;
        RECT 20.890 8.890 21.290 9.290 ;
        RECT 22.890 8.890 23.290 9.290 ;
        RECT 24.890 8.890 25.290 9.290 ;
        RECT 26.890 8.890 27.290 9.290 ;
        RECT 28.890 8.890 29.290 9.290 ;
        RECT 30.890 8.890 31.290 9.290 ;
        RECT 32.890 8.890 33.290 9.290 ;
        RECT 34.890 8.890 35.290 9.290 ;
        RECT 36.890 8.890 37.290 9.290 ;
        RECT 38.890 8.890 39.290 9.290 ;
        RECT 40.890 8.890 41.290 9.290 ;
        RECT 42.890 8.890 43.290 9.290 ;
        RECT 44.890 8.890 45.290 9.290 ;
        RECT 46.890 8.890 47.290 9.290 ;
        RECT 48.890 8.890 49.290 9.290 ;
        RECT 50.890 8.890 51.290 9.290 ;
        RECT 52.890 8.890 53.290 9.290 ;
        RECT 54.890 8.890 55.290 9.290 ;
        RECT 56.890 8.890 57.290 9.290 ;
        RECT 58.890 8.890 59.290 9.290 ;
        RECT 60.890 8.890 61.290 9.290 ;
        RECT 62.890 8.890 63.290 9.290 ;
        RECT 64.890 8.890 65.290 9.290 ;
        RECT 66.890 8.890 67.290 9.290 ;
        RECT 68.890 8.890 69.290 9.290 ;
        RECT 70.890 8.890 71.290 9.290 ;
        RECT 72.890 8.890 73.290 9.290 ;
        RECT 87.825 8.890 88.225 9.290 ;
        RECT 89.825 8.890 90.225 9.290 ;
        RECT 91.825 8.890 92.225 9.290 ;
        RECT 93.825 8.890 94.225 9.290 ;
        RECT 95.825 8.890 96.225 9.290 ;
        RECT 97.825 8.890 98.225 9.290 ;
        RECT 99.825 8.890 100.225 9.290 ;
        RECT 101.825 8.890 102.225 9.290 ;
        RECT 103.825 8.890 104.225 9.290 ;
        RECT 105.825 8.890 106.225 9.290 ;
        RECT 107.825 8.890 108.225 9.290 ;
        RECT 109.825 8.890 110.225 9.290 ;
        RECT 111.825 8.890 112.225 9.290 ;
        RECT 113.825 8.890 114.225 9.290 ;
        RECT 115.825 8.890 116.225 9.290 ;
        RECT 117.825 8.890 118.225 9.290 ;
        RECT 119.825 8.890 120.225 9.290 ;
        RECT 121.825 8.890 122.225 9.290 ;
        RECT 123.825 8.890 124.225 9.290 ;
        RECT 125.825 8.890 126.225 9.290 ;
        RECT 127.825 8.890 128.225 9.290 ;
        RECT 129.825 8.890 130.225 9.290 ;
        RECT 131.825 8.890 132.225 9.290 ;
        RECT 133.825 8.890 134.225 9.290 ;
        RECT 135.825 8.890 136.225 9.290 ;
        RECT 137.825 8.890 138.225 9.290 ;
        RECT 139.825 8.890 140.225 9.290 ;
        RECT 141.825 8.890 142.225 9.290 ;
        RECT 143.825 8.890 144.225 9.290 ;
        RECT 145.825 8.890 146.225 9.290 ;
        RECT 147.825 8.890 148.225 9.290 ;
        RECT 149.825 8.890 150.225 9.290 ;
        RECT 151.825 8.890 152.225 9.290 ;
        RECT 153.825 8.890 154.225 9.290 ;
        RECT 6.960 8.040 7.220 8.890 ;
        RECT 8.990 8.040 9.190 8.890 ;
        RECT 10.990 8.040 11.190 8.890 ;
        RECT 12.990 8.040 13.190 8.890 ;
        RECT 14.990 8.040 15.190 8.890 ;
        RECT 16.990 8.040 17.190 8.890 ;
        RECT 18.990 8.040 19.190 8.890 ;
        RECT 20.990 8.040 21.190 8.890 ;
        RECT 22.990 8.040 23.190 8.890 ;
        RECT 24.990 8.040 25.190 8.890 ;
        RECT 26.990 8.040 27.190 8.890 ;
        RECT 28.990 8.040 29.190 8.890 ;
        RECT 30.990 8.040 31.190 8.890 ;
        RECT 32.990 8.040 33.190 8.890 ;
        RECT 34.990 8.040 35.190 8.890 ;
        RECT 36.990 8.040 37.190 8.890 ;
        RECT 38.990 8.040 39.190 8.890 ;
        RECT 40.990 8.040 41.190 8.890 ;
        RECT 42.990 8.040 43.190 8.890 ;
        RECT 44.990 8.040 45.190 8.890 ;
        RECT 46.990 8.040 47.190 8.890 ;
        RECT 48.990 8.040 49.190 8.890 ;
        RECT 50.990 8.040 51.190 8.890 ;
        RECT 52.990 8.040 53.190 8.890 ;
        RECT 54.990 8.040 55.190 8.890 ;
        RECT 56.990 8.040 57.190 8.890 ;
        RECT 58.990 8.040 59.190 8.890 ;
        RECT 60.990 8.040 61.190 8.890 ;
        RECT 62.990 8.040 63.190 8.890 ;
        RECT 64.990 8.040 65.190 8.890 ;
        RECT 66.990 8.040 67.190 8.890 ;
        RECT 68.990 8.040 69.190 8.890 ;
        RECT 70.990 8.040 71.190 8.890 ;
        RECT 89.925 8.040 90.125 8.890 ;
        RECT 91.925 8.040 92.125 8.890 ;
        RECT 93.925 8.040 94.125 8.890 ;
        RECT 95.925 8.040 96.125 8.890 ;
        RECT 97.925 8.040 98.125 8.890 ;
        RECT 99.925 8.040 100.125 8.890 ;
        RECT 101.925 8.040 102.125 8.890 ;
        RECT 103.925 8.040 104.125 8.890 ;
        RECT 105.925 8.040 106.125 8.890 ;
        RECT 107.925 8.040 108.125 8.890 ;
        RECT 109.925 8.040 110.125 8.890 ;
        RECT 111.925 8.040 112.125 8.890 ;
        RECT 113.925 8.040 114.125 8.890 ;
        RECT 115.925 8.040 116.125 8.890 ;
        RECT 117.925 8.040 118.125 8.890 ;
        RECT 119.925 8.040 120.125 8.890 ;
        RECT 121.925 8.040 122.125 8.890 ;
        RECT 123.925 8.040 124.125 8.890 ;
        RECT 125.925 8.040 126.125 8.890 ;
        RECT 127.925 8.040 128.125 8.890 ;
        RECT 129.925 8.040 130.125 8.890 ;
        RECT 131.925 8.040 132.125 8.890 ;
        RECT 133.925 8.040 134.125 8.890 ;
        RECT 135.925 8.040 136.125 8.890 ;
        RECT 137.925 8.040 138.125 8.890 ;
        RECT 139.925 8.040 140.125 8.890 ;
        RECT 141.925 8.040 142.125 8.890 ;
        RECT 143.925 8.040 144.125 8.890 ;
        RECT 145.925 8.040 146.125 8.890 ;
        RECT 147.925 8.040 148.125 8.890 ;
        RECT 149.925 8.040 150.125 8.890 ;
        RECT 151.925 8.040 152.125 8.890 ;
        RECT 153.895 8.040 154.155 8.890 ;
        RECT 6.890 7.640 7.290 8.040 ;
        RECT 8.890 7.640 9.290 8.040 ;
        RECT 10.890 7.640 11.290 8.040 ;
        RECT 12.890 7.640 13.290 8.040 ;
        RECT 14.890 7.640 15.290 8.040 ;
        RECT 16.890 7.640 17.290 8.040 ;
        RECT 18.890 7.640 19.290 8.040 ;
        RECT 20.890 7.640 21.290 8.040 ;
        RECT 22.890 7.640 23.290 8.040 ;
        RECT 24.890 7.640 25.290 8.040 ;
        RECT 26.890 7.640 27.290 8.040 ;
        RECT 28.890 7.640 29.290 8.040 ;
        RECT 30.890 7.640 31.290 8.040 ;
        RECT 32.890 7.640 33.290 8.040 ;
        RECT 34.890 7.640 35.290 8.040 ;
        RECT 36.890 7.640 37.290 8.040 ;
        RECT 38.890 7.640 39.290 8.040 ;
        RECT 40.890 7.640 41.290 8.040 ;
        RECT 42.890 7.640 43.290 8.040 ;
        RECT 44.890 7.640 45.290 8.040 ;
        RECT 46.890 7.640 47.290 8.040 ;
        RECT 48.890 7.640 49.290 8.040 ;
        RECT 50.890 7.640 51.290 8.040 ;
        RECT 52.890 7.640 53.290 8.040 ;
        RECT 54.890 7.640 55.290 8.040 ;
        RECT 56.890 7.640 57.290 8.040 ;
        RECT 58.890 7.640 59.290 8.040 ;
        RECT 60.890 7.640 61.290 8.040 ;
        RECT 62.890 7.640 63.290 8.040 ;
        RECT 64.890 7.640 65.290 8.040 ;
        RECT 66.890 7.640 67.290 8.040 ;
        RECT 68.890 7.640 69.290 8.040 ;
        RECT 70.890 7.640 71.290 8.040 ;
        RECT 72.890 7.640 73.290 8.040 ;
        RECT 87.825 7.640 88.225 8.040 ;
        RECT 89.825 7.640 90.225 8.040 ;
        RECT 91.825 7.640 92.225 8.040 ;
        RECT 93.825 7.640 94.225 8.040 ;
        RECT 95.825 7.640 96.225 8.040 ;
        RECT 97.825 7.640 98.225 8.040 ;
        RECT 99.825 7.640 100.225 8.040 ;
        RECT 101.825 7.640 102.225 8.040 ;
        RECT 103.825 7.640 104.225 8.040 ;
        RECT 105.825 7.640 106.225 8.040 ;
        RECT 107.825 7.640 108.225 8.040 ;
        RECT 109.825 7.640 110.225 8.040 ;
        RECT 111.825 7.640 112.225 8.040 ;
        RECT 113.825 7.640 114.225 8.040 ;
        RECT 115.825 7.640 116.225 8.040 ;
        RECT 117.825 7.640 118.225 8.040 ;
        RECT 119.825 7.640 120.225 8.040 ;
        RECT 121.825 7.640 122.225 8.040 ;
        RECT 123.825 7.640 124.225 8.040 ;
        RECT 125.825 7.640 126.225 8.040 ;
        RECT 127.825 7.640 128.225 8.040 ;
        RECT 129.825 7.640 130.225 8.040 ;
        RECT 131.825 7.640 132.225 8.040 ;
        RECT 133.825 7.640 134.225 8.040 ;
        RECT 135.825 7.640 136.225 8.040 ;
        RECT 137.825 7.640 138.225 8.040 ;
        RECT 139.825 7.640 140.225 8.040 ;
        RECT 141.825 7.640 142.225 8.040 ;
        RECT 143.825 7.640 144.225 8.040 ;
        RECT 145.825 7.640 146.225 8.040 ;
        RECT 147.825 7.640 148.225 8.040 ;
        RECT 149.825 7.640 150.225 8.040 ;
        RECT 151.825 7.640 152.225 8.040 ;
        RECT 153.825 7.640 154.225 8.040 ;
        RECT 6.890 7.440 8.540 7.640 ;
        RECT 8.890 7.440 74.540 7.640 ;
        RECT 86.575 7.440 152.225 7.640 ;
        RECT 152.575 7.440 154.225 7.640 ;
        RECT 6.890 7.040 7.290 7.440 ;
        RECT 8.890 7.040 9.290 7.440 ;
        RECT 10.890 7.040 11.290 7.440 ;
        RECT 12.890 7.040 13.290 7.440 ;
        RECT 14.890 7.040 15.290 7.440 ;
        RECT 16.890 7.040 17.290 7.440 ;
        RECT 18.890 7.040 19.290 7.440 ;
        RECT 20.890 7.040 21.290 7.440 ;
        RECT 22.890 7.040 23.290 7.440 ;
        RECT 24.890 7.040 25.290 7.440 ;
        RECT 26.890 7.040 27.290 7.440 ;
        RECT 28.890 7.040 29.290 7.440 ;
        RECT 30.890 7.040 31.290 7.440 ;
        RECT 32.890 7.040 33.290 7.440 ;
        RECT 34.890 7.040 35.290 7.440 ;
        RECT 36.890 7.040 37.290 7.440 ;
        RECT 38.890 7.040 39.290 7.440 ;
        RECT 40.890 7.040 41.290 7.440 ;
        RECT 42.890 7.040 43.290 7.440 ;
        RECT 44.890 7.040 45.290 7.440 ;
        RECT 46.890 7.040 47.290 7.440 ;
        RECT 48.890 7.040 49.290 7.440 ;
        RECT 50.890 7.040 51.290 7.440 ;
        RECT 52.890 7.040 53.290 7.440 ;
        RECT 54.890 7.040 55.290 7.440 ;
        RECT 56.890 7.040 57.290 7.440 ;
        RECT 58.890 7.040 59.290 7.440 ;
        RECT 60.890 7.040 61.290 7.440 ;
        RECT 62.890 7.040 63.290 7.440 ;
        RECT 64.890 7.040 65.290 7.440 ;
        RECT 66.890 7.040 67.290 7.440 ;
        RECT 68.890 7.040 69.290 7.440 ;
        RECT 70.890 7.040 71.290 7.440 ;
        RECT 72.890 7.040 73.290 7.440 ;
        RECT 87.825 7.040 88.225 7.440 ;
        RECT 89.825 7.040 90.225 7.440 ;
        RECT 91.825 7.040 92.225 7.440 ;
        RECT 93.825 7.040 94.225 7.440 ;
        RECT 95.825 7.040 96.225 7.440 ;
        RECT 97.825 7.040 98.225 7.440 ;
        RECT 99.825 7.040 100.225 7.440 ;
        RECT 101.825 7.040 102.225 7.440 ;
        RECT 103.825 7.040 104.225 7.440 ;
        RECT 105.825 7.040 106.225 7.440 ;
        RECT 107.825 7.040 108.225 7.440 ;
        RECT 109.825 7.040 110.225 7.440 ;
        RECT 111.825 7.040 112.225 7.440 ;
        RECT 113.825 7.040 114.225 7.440 ;
        RECT 115.825 7.040 116.225 7.440 ;
        RECT 117.825 7.040 118.225 7.440 ;
        RECT 119.825 7.040 120.225 7.440 ;
        RECT 121.825 7.040 122.225 7.440 ;
        RECT 123.825 7.040 124.225 7.440 ;
        RECT 125.825 7.040 126.225 7.440 ;
        RECT 127.825 7.040 128.225 7.440 ;
        RECT 129.825 7.040 130.225 7.440 ;
        RECT 131.825 7.040 132.225 7.440 ;
        RECT 133.825 7.040 134.225 7.440 ;
        RECT 135.825 7.040 136.225 7.440 ;
        RECT 137.825 7.040 138.225 7.440 ;
        RECT 139.825 7.040 140.225 7.440 ;
        RECT 141.825 7.040 142.225 7.440 ;
        RECT 143.825 7.040 144.225 7.440 ;
        RECT 145.825 7.040 146.225 7.440 ;
        RECT 147.825 7.040 148.225 7.440 ;
        RECT 149.825 7.040 150.225 7.440 ;
        RECT 151.825 7.040 152.225 7.440 ;
        RECT 153.825 7.040 154.225 7.440 ;
        RECT 6.960 6.190 7.220 7.040 ;
        RECT 153.895 6.190 154.155 7.040 ;
        RECT 6.890 5.790 7.290 6.190 ;
        RECT 8.890 5.820 9.290 6.190 ;
        RECT 10.890 5.820 11.290 6.190 ;
        RECT 12.890 5.820 13.290 6.190 ;
        RECT 14.890 5.820 15.290 6.190 ;
        RECT 16.890 5.820 17.290 6.190 ;
        RECT 18.890 5.820 19.290 6.190 ;
        RECT 20.890 5.820 21.290 6.190 ;
        RECT 22.890 5.820 23.290 6.190 ;
        RECT 24.890 5.820 25.290 6.190 ;
        RECT 26.890 5.820 27.290 6.190 ;
        RECT 28.890 5.820 29.290 6.190 ;
        RECT 30.890 5.820 31.290 6.190 ;
        RECT 32.890 5.820 33.290 6.190 ;
        RECT 34.890 5.820 35.290 6.190 ;
        RECT 36.890 5.820 37.290 6.190 ;
        RECT 38.890 5.820 39.290 6.190 ;
        RECT 40.890 5.820 41.290 6.190 ;
        RECT 42.890 5.820 43.290 6.190 ;
        RECT 44.890 5.820 45.290 6.190 ;
        RECT 46.890 5.820 47.290 6.190 ;
        RECT 48.890 5.820 49.290 6.190 ;
        RECT 50.890 5.820 51.290 6.190 ;
        RECT 52.890 5.820 53.290 6.190 ;
        RECT 54.890 5.820 55.290 6.190 ;
        RECT 56.890 5.820 57.290 6.190 ;
        RECT 58.890 5.820 59.290 6.190 ;
        RECT 60.890 5.820 61.290 6.190 ;
        RECT 62.890 5.820 63.290 6.190 ;
        RECT 64.890 5.820 65.290 6.190 ;
        RECT 66.890 5.820 67.290 6.190 ;
        RECT 68.890 5.820 69.290 6.190 ;
        RECT 70.890 5.820 71.290 6.190 ;
        RECT 72.890 5.820 73.290 6.190 ;
        RECT 87.825 5.820 88.225 6.190 ;
        RECT 89.825 5.820 90.225 6.190 ;
        RECT 91.825 5.820 92.225 6.190 ;
        RECT 93.825 5.820 94.225 6.190 ;
        RECT 95.825 5.820 96.225 6.190 ;
        RECT 97.825 5.820 98.225 6.190 ;
        RECT 99.825 5.820 100.225 6.190 ;
        RECT 101.825 5.820 102.225 6.190 ;
        RECT 103.825 5.820 104.225 6.190 ;
        RECT 105.825 5.820 106.225 6.190 ;
        RECT 107.825 5.820 108.225 6.190 ;
        RECT 109.825 5.820 110.225 6.190 ;
        RECT 111.825 5.820 112.225 6.190 ;
        RECT 113.825 5.820 114.225 6.190 ;
        RECT 115.825 5.820 116.225 6.190 ;
        RECT 117.825 5.820 118.225 6.190 ;
        RECT 119.825 5.820 120.225 6.190 ;
        RECT 121.825 5.820 122.225 6.190 ;
        RECT 123.825 5.820 124.225 6.190 ;
        RECT 125.825 5.820 126.225 6.190 ;
        RECT 127.825 5.820 128.225 6.190 ;
        RECT 129.825 5.820 130.225 6.190 ;
        RECT 131.825 5.820 132.225 6.190 ;
        RECT 133.825 5.820 134.225 6.190 ;
        RECT 135.825 5.820 136.225 6.190 ;
        RECT 137.825 5.820 138.225 6.190 ;
        RECT 139.825 5.820 140.225 6.190 ;
        RECT 141.825 5.820 142.225 6.190 ;
        RECT 143.825 5.820 144.225 6.190 ;
        RECT 145.825 5.820 146.225 6.190 ;
        RECT 147.825 5.820 148.225 6.190 ;
        RECT 149.825 5.820 150.225 6.190 ;
        RECT 151.825 5.820 152.225 6.190 ;
        RECT 7.680 5.790 73.700 5.820 ;
        RECT 87.415 5.790 153.435 5.820 ;
        RECT 153.825 5.790 154.225 6.190 ;
        RECT 6.890 5.590 74.540 5.790 ;
        RECT 86.575 5.590 154.225 5.790 ;
        RECT 6.890 5.190 7.290 5.590 ;
        RECT 7.680 5.560 73.700 5.590 ;
        RECT 87.415 5.560 153.435 5.590 ;
        RECT 8.890 5.190 9.290 5.560 ;
        RECT 10.890 5.190 11.290 5.560 ;
        RECT 12.890 5.190 13.290 5.560 ;
        RECT 14.890 5.190 15.290 5.560 ;
        RECT 16.890 5.190 17.290 5.560 ;
        RECT 18.890 5.190 19.290 5.560 ;
        RECT 20.890 5.190 21.290 5.560 ;
        RECT 22.890 5.190 23.290 5.560 ;
        RECT 24.890 5.190 25.290 5.560 ;
        RECT 26.890 5.190 27.290 5.560 ;
        RECT 28.890 5.190 29.290 5.560 ;
        RECT 30.890 5.190 31.290 5.560 ;
        RECT 32.890 5.190 33.290 5.560 ;
        RECT 34.890 5.190 35.290 5.560 ;
        RECT 36.890 5.190 37.290 5.560 ;
        RECT 38.890 5.190 39.290 5.560 ;
        RECT 40.890 5.190 41.290 5.560 ;
        RECT 42.890 5.190 43.290 5.560 ;
        RECT 44.890 5.190 45.290 5.560 ;
        RECT 46.890 5.190 47.290 5.560 ;
        RECT 48.890 5.190 49.290 5.560 ;
        RECT 50.890 5.190 51.290 5.560 ;
        RECT 52.890 5.190 53.290 5.560 ;
        RECT 54.890 5.190 55.290 5.560 ;
        RECT 56.890 5.190 57.290 5.560 ;
        RECT 58.890 5.190 59.290 5.560 ;
        RECT 60.890 5.190 61.290 5.560 ;
        RECT 62.890 5.190 63.290 5.560 ;
        RECT 64.890 5.190 65.290 5.560 ;
        RECT 66.890 5.190 67.290 5.560 ;
        RECT 68.890 5.190 69.290 5.560 ;
        RECT 70.890 5.190 71.290 5.560 ;
        RECT 72.890 5.190 73.290 5.560 ;
        RECT 87.825 5.190 88.225 5.560 ;
        RECT 89.825 5.190 90.225 5.560 ;
        RECT 91.825 5.190 92.225 5.560 ;
        RECT 93.825 5.190 94.225 5.560 ;
        RECT 95.825 5.190 96.225 5.560 ;
        RECT 97.825 5.190 98.225 5.560 ;
        RECT 99.825 5.190 100.225 5.560 ;
        RECT 101.825 5.190 102.225 5.560 ;
        RECT 103.825 5.190 104.225 5.560 ;
        RECT 105.825 5.190 106.225 5.560 ;
        RECT 107.825 5.190 108.225 5.560 ;
        RECT 109.825 5.190 110.225 5.560 ;
        RECT 111.825 5.190 112.225 5.560 ;
        RECT 113.825 5.190 114.225 5.560 ;
        RECT 115.825 5.190 116.225 5.560 ;
        RECT 117.825 5.190 118.225 5.560 ;
        RECT 119.825 5.190 120.225 5.560 ;
        RECT 121.825 5.190 122.225 5.560 ;
        RECT 123.825 5.190 124.225 5.560 ;
        RECT 125.825 5.190 126.225 5.560 ;
        RECT 127.825 5.190 128.225 5.560 ;
        RECT 129.825 5.190 130.225 5.560 ;
        RECT 131.825 5.190 132.225 5.560 ;
        RECT 133.825 5.190 134.225 5.560 ;
        RECT 135.825 5.190 136.225 5.560 ;
        RECT 137.825 5.190 138.225 5.560 ;
        RECT 139.825 5.190 140.225 5.560 ;
        RECT 141.825 5.190 142.225 5.560 ;
        RECT 143.825 5.190 144.225 5.560 ;
        RECT 145.825 5.190 146.225 5.560 ;
        RECT 147.825 5.190 148.225 5.560 ;
        RECT 149.825 5.190 150.225 5.560 ;
        RECT 151.825 5.190 152.225 5.560 ;
        RECT 153.825 5.190 154.225 5.590 ;
      LAYER met2 ;
        RECT 14.850 223.075 15.150 223.475 ;
        RECT 10.215 219.490 10.515 219.640 ;
        RECT 12.140 219.490 12.440 219.690 ;
        RECT 10.215 219.340 12.440 219.490 ;
        RECT 10.215 219.240 10.515 219.340 ;
        RECT 12.140 219.290 12.440 219.340 ;
        RECT 14.410 219.310 14.690 219.680 ;
        RECT 14.480 218.465 14.620 219.310 ;
        RECT 9.815 218.190 10.115 218.340 ;
        RECT 12.140 218.190 12.440 218.290 ;
        RECT 9.815 218.040 12.440 218.190 ;
        RECT 9.815 217.940 10.115 218.040 ;
        RECT 12.140 217.890 12.440 218.040 ;
        RECT 13.950 217.950 14.230 218.320 ;
        RECT 14.420 218.145 14.680 218.465 ;
        RECT 14.870 218.265 15.150 223.075 ;
        RECT 134.450 223.050 134.750 223.450 ;
        RECT 26.810 222.425 27.110 222.825 ;
        RECT 14.020 217.445 14.160 217.950 ;
        RECT 13.960 217.125 14.220 217.445 ;
        RECT 14.940 217.105 15.080 218.265 ;
        RECT 21.780 218.145 22.040 218.465 ;
        RECT 22.700 218.145 22.960 218.465 ;
        RECT 26.830 218.265 27.110 222.425 ;
        RECT 38.770 221.825 39.070 222.225 ;
        RECT 122.500 221.900 122.800 222.300 ;
        RECT 38.790 218.265 39.070 221.825 ;
        RECT 50.730 221.225 51.040 221.625 ;
        RECT 98.600 221.590 98.900 221.650 ;
        RECT 45.700 219.165 45.960 219.485 ;
        RECT 50.750 219.340 51.040 221.225 ;
        RECT 98.590 221.250 98.900 221.590 ;
        RECT 62.690 220.625 62.990 221.025 ;
        RECT 43.400 218.485 43.660 218.805 ;
        RECT 9.465 216.840 9.765 216.990 ;
        RECT 12.140 216.840 12.440 216.990 ;
        RECT 9.465 216.690 12.440 216.840 ;
        RECT 14.880 216.785 15.140 217.105 ;
        RECT 9.465 216.590 9.765 216.690 ;
        RECT 12.140 216.590 12.440 216.690 ;
        RECT 17.630 216.590 17.910 216.960 ;
        RECT 21.310 216.590 21.590 216.960 ;
        RECT 21.840 216.765 21.980 218.145 ;
        RECT 22.760 217.445 22.900 218.145 ;
        RECT 22.700 217.125 22.960 217.445 ;
        RECT 22.240 216.785 22.500 217.105 ;
        RECT 9.165 215.440 9.465 215.590 ;
        RECT 12.140 215.440 12.440 215.590 ;
        RECT 9.165 215.290 12.440 215.440 ;
        RECT 9.165 215.190 9.465 215.290 ;
        RECT 12.140 215.190 12.440 215.290 ;
        RECT 15.790 215.230 16.070 215.600 ;
        RECT 15.860 214.725 16.000 215.230 ;
        RECT 17.700 214.725 17.840 216.590 ;
        RECT 21.320 216.445 21.580 216.590 ;
        RECT 21.780 216.445 22.040 216.765 ;
        RECT 20.400 215.425 20.660 215.745 ;
        RECT 15.800 214.405 16.060 214.725 ;
        RECT 17.640 214.405 17.900 214.725 ;
        RECT 20.460 214.240 20.600 215.425 ;
        RECT 21.780 214.240 22.040 214.385 ;
        RECT 8.865 214.090 9.165 214.240 ;
        RECT 12.090 214.090 12.390 214.240 ;
        RECT 8.865 213.940 12.390 214.090 ;
        RECT 8.865 213.840 9.165 213.940 ;
        RECT 12.090 213.840 12.390 213.940 ;
        RECT 19.020 213.725 19.280 214.045 ;
        RECT 20.390 213.870 20.670 214.240 ;
        RECT 21.770 213.870 22.050 214.240 ;
        RECT 8.565 212.690 8.865 212.840 ;
        RECT 12.090 212.690 12.390 212.890 ;
        RECT 14.420 212.705 14.680 213.025 ;
        RECT 8.565 212.540 12.390 212.690 ;
        RECT 8.565 212.440 8.865 212.540 ;
        RECT 12.090 212.490 12.390 212.540 ;
        RECT 8.265 211.390 8.565 211.540 ;
        RECT 12.140 211.390 12.440 211.540 ;
        RECT 14.480 211.520 14.620 212.705 ;
        RECT 14.870 212.510 15.150 212.880 ;
        RECT 14.940 212.005 15.080 212.510 ;
        RECT 14.880 211.685 15.140 212.005 ;
        RECT 8.265 211.240 12.440 211.390 ;
        RECT 8.265 211.140 8.565 211.240 ;
        RECT 12.140 211.140 12.440 211.240 ;
        RECT 14.410 211.150 14.690 211.520 ;
        RECT 19.080 211.325 19.220 213.725 ;
        RECT 19.480 213.385 19.740 213.705 ;
        RECT 20.400 213.560 20.660 213.705 ;
        RECT 18.560 211.005 18.820 211.325 ;
        RECT 19.020 211.005 19.280 211.325 ;
        RECT 14.540 210.325 14.800 210.645 ;
        RECT 7.965 210.040 8.265 210.190 ;
        RECT 12.090 210.040 12.390 210.190 ;
        RECT 14.600 210.160 14.740 210.325 ;
        RECT 7.965 209.890 12.390 210.040 ;
        RECT 7.965 209.790 8.265 209.890 ;
        RECT 12.090 209.790 12.390 209.890 ;
        RECT 14.530 209.790 14.810 210.160 ;
        RECT 7.665 208.640 7.965 208.790 ;
        RECT 12.140 208.640 12.440 208.840 ;
        RECT 14.200 208.800 14.460 208.945 ;
        RECT 18.620 208.800 18.760 211.005 ;
        RECT 7.665 208.490 12.440 208.640 ;
        RECT 7.665 208.390 7.965 208.490 ;
        RECT 12.140 208.440 12.440 208.490 ;
        RECT 14.190 208.430 14.470 208.800 ;
        RECT 18.550 208.430 18.830 208.800 ;
        RECT 16.720 208.120 16.980 208.265 ;
        RECT 16.710 207.750 16.990 208.120 ;
        RECT 7.365 207.290 7.665 207.440 ;
        RECT 12.140 207.290 12.440 207.490 ;
        RECT 17.640 207.440 17.900 207.585 ;
        RECT 7.365 207.140 12.440 207.290 ;
        RECT 7.365 207.040 7.665 207.140 ;
        RECT 12.140 207.090 12.440 207.140 ;
        RECT 17.630 207.070 17.910 207.440 ;
        RECT 14.120 206.245 14.380 206.565 ;
        RECT 7.065 205.990 7.365 206.140 ;
        RECT 12.140 205.990 12.440 206.090 ;
        RECT 14.180 206.080 14.320 206.245 ;
        RECT 7.065 205.840 12.440 205.990 ;
        RECT 7.065 205.740 7.365 205.840 ;
        RECT 12.140 205.690 12.440 205.840 ;
        RECT 14.110 205.710 14.390 206.080 ;
        RECT 17.170 205.030 17.450 205.400 ;
        RECT 6.765 204.590 7.065 204.740 ;
        RECT 12.140 204.590 12.440 204.740 ;
        RECT 14.090 204.720 14.350 204.865 ;
        RECT 6.765 204.440 12.440 204.590 ;
        RECT 6.765 204.340 7.065 204.440 ;
        RECT 12.140 204.340 12.440 204.440 ;
        RECT 14.080 204.350 14.360 204.720 ;
        RECT 6.465 203.240 6.765 203.390 ;
        RECT 13.960 203.360 14.220 203.505 ;
        RECT 12.140 203.240 12.440 203.340 ;
        RECT 6.465 203.090 12.440 203.240 ;
        RECT 6.465 202.990 6.765 203.090 ;
        RECT 12.140 202.940 12.440 203.090 ;
        RECT 13.950 202.990 14.230 203.360 ;
        RECT 16.710 202.990 16.990 203.360 ;
        RECT 16.780 202.825 16.920 202.990 ;
        RECT 16.720 202.505 16.980 202.825 ;
        RECT 6.165 201.840 6.465 201.990 ;
        RECT 12.140 201.840 12.440 201.990 ;
        RECT 6.165 201.690 12.440 201.840 ;
        RECT 6.165 201.590 6.465 201.690 ;
        RECT 12.140 201.590 12.440 201.690 ;
        RECT 15.790 201.630 16.070 202.000 ;
        RECT 5.865 200.540 6.165 200.690 ;
        RECT 12.140 200.540 12.440 200.640 ;
        RECT 5.865 200.390 12.440 200.540 ;
        RECT 5.865 200.290 6.165 200.390 ;
        RECT 12.140 200.240 12.440 200.390 ;
        RECT 15.860 199.765 16.000 201.630 ;
        RECT 15.800 199.445 16.060 199.765 ;
        RECT 16.710 199.590 16.990 199.960 ;
        RECT 5.565 199.190 5.865 199.340 ;
        RECT 12.140 199.190 12.440 199.290 ;
        RECT 5.565 199.040 12.440 199.190 ;
        RECT 5.565 198.940 5.865 199.040 ;
        RECT 12.140 198.890 12.440 199.040 ;
        RECT 14.870 198.910 15.150 199.280 ;
        RECT 14.940 198.405 15.080 198.910 ;
        RECT 14.880 198.085 15.140 198.405 ;
        RECT 5.265 197.840 5.565 197.990 ;
        RECT 12.140 197.840 12.440 197.940 ;
        RECT 5.265 197.690 12.440 197.840 ;
        RECT 5.265 197.590 5.565 197.690 ;
        RECT 12.140 197.540 12.440 197.690 ;
        RECT 14.410 197.550 14.690 197.920 ;
        RECT 4.965 196.390 5.265 196.540 ;
        RECT 12.140 196.390 12.440 196.590 ;
        RECT 4.965 196.240 12.440 196.390 ;
        RECT 4.965 196.140 5.265 196.240 ;
        RECT 12.140 196.190 12.440 196.240 ;
        RECT 4.665 195.040 4.965 195.190 ;
        RECT 12.140 195.040 12.440 195.240 ;
        RECT 4.665 194.890 12.440 195.040 ;
        RECT 4.665 194.790 4.965 194.890 ;
        RECT 12.140 194.840 12.440 194.890 ;
        RECT 14.480 194.325 14.620 197.550 ;
        RECT 14.870 196.190 15.150 196.560 ;
        RECT 14.940 195.685 15.080 196.190 ;
        RECT 14.880 195.365 15.140 195.685 ;
        RECT 15.790 194.830 16.070 195.200 ;
        RECT 16.780 195.005 16.920 199.590 ;
        RECT 17.240 197.385 17.380 205.030 ;
        RECT 18.560 204.545 18.820 204.865 ;
        RECT 18.090 202.310 18.370 202.680 ;
        RECT 17.630 200.270 17.910 200.640 ;
        RECT 18.160 200.445 18.300 202.310 ;
        RECT 17.700 199.765 17.840 200.270 ;
        RECT 18.100 200.125 18.360 200.445 ;
        RECT 17.640 199.445 17.900 199.765 ;
        RECT 17.180 197.065 17.440 197.385 ;
        RECT 14.420 194.005 14.680 194.325 ;
        RECT 4.365 193.740 4.665 193.890 ;
        RECT 12.140 193.740 12.440 193.890 ;
        RECT 4.365 193.590 12.440 193.740 ;
        RECT 4.365 193.490 4.665 193.590 ;
        RECT 12.140 193.490 12.440 193.590 ;
        RECT 15.860 192.965 16.000 194.830 ;
        RECT 16.720 194.685 16.980 195.005 ;
        RECT 18.090 194.830 18.370 195.200 ;
        RECT 18.100 194.685 18.360 194.830 ;
        RECT 17.630 193.470 17.910 193.840 ;
        RECT 17.700 192.965 17.840 193.470 ;
        RECT 15.800 192.645 16.060 192.965 ;
        RECT 17.640 192.645 17.900 192.965 ;
        RECT 4.065 192.290 4.365 192.440 ;
        RECT 12.140 192.290 12.440 192.540 ;
        RECT 4.065 192.140 12.440 192.290 ;
        RECT 4.065 192.040 4.365 192.140 ;
        RECT 13.490 192.110 13.770 192.480 ;
        RECT 14.880 192.305 15.140 192.625 ;
        RECT 13.560 191.265 13.700 192.110 ;
        RECT 13.960 191.965 14.220 192.285 ;
        RECT 3.765 190.940 4.065 191.090 ;
        RECT 12.140 190.940 12.440 191.190 ;
        RECT 13.500 190.945 13.760 191.265 ;
        RECT 3.765 190.790 12.440 190.940 ;
        RECT 3.765 190.690 4.065 190.790 ;
        RECT 3.465 189.540 3.765 189.690 ;
        RECT 12.140 189.540 12.440 189.640 ;
        RECT 3.465 189.390 12.440 189.540 ;
        RECT 3.465 189.290 3.765 189.390 ;
        RECT 12.140 189.240 12.440 189.390 ;
        RECT 14.020 187.715 14.160 191.965 ;
        RECT 14.940 191.120 15.080 192.305 ;
        RECT 16.720 191.625 16.980 191.945 ;
        RECT 14.870 190.750 15.150 191.120 ;
        RECT 16.780 189.905 16.920 191.625 ;
        RECT 16.720 189.585 16.980 189.905 ;
        RECT 18.620 187.715 18.760 204.545 ;
        RECT 19.080 203.165 19.220 211.005 ;
        RECT 19.540 206.080 19.680 213.385 ;
        RECT 20.390 213.190 20.670 213.560 ;
        RECT 19.470 205.710 19.750 206.080 ;
        RECT 19.940 205.565 20.200 205.885 ;
        RECT 19.020 202.845 19.280 203.165 ;
        RECT 19.080 200.445 19.220 202.845 ;
        RECT 19.020 200.125 19.280 200.445 ;
        RECT 19.080 197.725 19.220 200.125 ;
        RECT 19.480 199.445 19.740 199.765 ;
        RECT 19.020 197.405 19.280 197.725 ;
        RECT 19.080 195.005 19.220 197.405 ;
        RECT 19.020 194.685 19.280 195.005 ;
        RECT 19.540 188.875 19.680 199.445 ;
        RECT 20.000 192.480 20.140 205.565 ;
        RECT 21.780 204.885 22.040 205.205 ;
        RECT 21.840 203.165 21.980 204.885 ;
        RECT 21.780 202.845 22.040 203.165 ;
        RECT 22.300 197.725 22.440 216.785 ;
        RECT 24.990 215.910 25.270 216.280 ;
        RECT 25.060 213.705 25.200 215.910 ;
        RECT 26.900 215.745 27.040 218.265 ;
        RECT 32.710 217.610 34.250 217.980 ;
        RECT 38.860 217.445 39.000 218.265 ;
        RECT 38.800 217.125 39.060 217.445 ;
        RECT 40.630 217.270 40.910 217.640 ;
        RECT 39.260 216.785 39.520 217.105 ;
        RECT 31.440 216.445 31.700 216.765 ;
        RECT 31.900 216.445 32.160 216.765 ;
        RECT 30.060 216.335 30.320 216.425 ;
        RECT 28.740 216.195 30.320 216.335 ;
        RECT 26.840 215.425 27.100 215.745 ;
        RECT 25.000 213.385 25.260 213.705 ;
        RECT 25.460 213.385 25.720 213.705 ;
        RECT 22.700 207.945 22.960 208.265 ;
        RECT 24.540 207.945 24.800 208.265 ;
        RECT 22.760 205.205 22.900 207.945 ;
        RECT 24.080 205.225 24.340 205.545 ;
        RECT 22.700 204.885 22.960 205.205 ;
        RECT 24.140 199.425 24.280 205.225 ;
        RECT 24.080 199.105 24.340 199.425 ;
        RECT 24.600 198.600 24.740 207.945 ;
        RECT 25.060 207.495 25.200 213.385 ;
        RECT 25.520 211.520 25.660 213.385 ;
        RECT 25.450 211.150 25.730 211.520 ;
        RECT 26.830 211.150 27.110 211.520 ;
        RECT 26.380 210.325 26.640 210.645 ;
        RECT 25.060 207.355 26.120 207.495 ;
        RECT 25.460 205.565 25.720 205.885 ;
        RECT 25.000 204.545 25.260 204.865 ;
        RECT 24.530 198.230 24.810 198.600 ;
        RECT 24.540 197.745 24.800 198.065 ;
        RECT 22.240 197.405 22.500 197.725 ;
        RECT 24.600 197.385 24.740 197.745 ;
        RECT 24.540 197.065 24.800 197.385 ;
        RECT 19.930 192.110 20.210 192.480 ;
        RECT 25.060 191.945 25.200 204.545 ;
        RECT 25.520 194.325 25.660 205.565 ;
        RECT 25.980 202.145 26.120 207.355 ;
        RECT 26.440 202.485 26.580 210.325 ;
        RECT 26.900 205.885 27.040 211.150 ;
        RECT 27.300 210.665 27.560 210.985 ;
        RECT 27.360 209.285 27.500 210.665 ;
        RECT 27.300 208.965 27.560 209.285 ;
        RECT 27.760 208.625 28.020 208.945 ;
        RECT 27.820 207.925 27.960 208.625 ;
        RECT 28.740 208.605 28.880 216.195 ;
        RECT 30.060 216.105 30.320 216.195 ;
        RECT 29.410 214.890 30.950 215.260 ;
        RECT 29.600 214.405 29.860 214.725 ;
        RECT 29.660 211.665 29.800 214.405 ;
        RECT 30.520 213.045 30.780 213.365 ;
        RECT 30.580 212.005 30.720 213.045 ;
        RECT 30.520 211.685 30.780 212.005 ;
        RECT 29.600 211.345 29.860 211.665 ;
        RECT 29.410 209.450 30.950 209.820 ;
        RECT 30.520 208.965 30.780 209.285 ;
        RECT 28.680 208.285 28.940 208.605 ;
        RECT 28.220 207.945 28.480 208.265 ;
        RECT 27.760 207.605 28.020 207.925 ;
        RECT 27.300 205.905 27.560 206.225 ;
        RECT 26.840 205.565 27.100 205.885 ;
        RECT 26.380 202.165 26.640 202.485 ;
        RECT 25.920 201.825 26.180 202.145 ;
        RECT 26.440 200.445 26.580 202.165 ;
        RECT 26.840 201.825 27.100 202.145 ;
        RECT 27.360 201.885 27.500 205.905 ;
        RECT 28.280 205.885 28.420 207.945 ;
        RECT 28.680 207.265 28.940 207.585 ;
        RECT 28.740 206.135 28.880 207.265 ;
        RECT 30.580 206.760 30.720 208.965 ;
        RECT 30.980 207.945 31.240 208.265 ;
        RECT 30.510 206.390 30.790 206.760 ;
        RECT 29.140 206.135 29.400 206.225 ;
        RECT 28.740 205.995 29.400 206.135 ;
        RECT 28.220 205.565 28.480 205.885 ;
        RECT 27.760 204.545 28.020 204.865 ;
        RECT 27.820 202.825 27.960 204.545 ;
        RECT 27.760 202.505 28.020 202.825 ;
        RECT 26.380 200.355 26.640 200.445 ;
        RECT 25.980 200.215 26.640 200.355 ;
        RECT 25.980 198.065 26.120 200.215 ;
        RECT 26.380 200.125 26.640 200.215 ;
        RECT 26.370 198.230 26.650 198.600 ;
        RECT 25.920 197.745 26.180 198.065 ;
        RECT 25.980 195.005 26.120 197.745 ;
        RECT 26.440 196.705 26.580 198.230 ;
        RECT 26.380 196.385 26.640 196.705 ;
        RECT 25.920 194.685 26.180 195.005 ;
        RECT 25.460 194.005 25.720 194.325 ;
        RECT 19.940 191.625 20.200 191.945 ;
        RECT 20.400 191.625 20.660 191.945 ;
        RECT 25.000 191.625 25.260 191.945 ;
        RECT 20.000 190.245 20.140 191.625 ;
        RECT 19.940 189.925 20.200 190.245 ;
        RECT 20.460 189.225 20.600 191.625 ;
        RECT 26.900 191.605 27.040 201.825 ;
        RECT 27.360 201.745 27.960 201.885 ;
        RECT 27.300 199.785 27.560 200.105 ;
        RECT 27.360 192.965 27.500 199.785 ;
        RECT 27.820 193.985 27.960 201.745 ;
        RECT 28.280 200.105 28.420 205.565 ;
        RECT 28.740 202.735 28.880 205.995 ;
        RECT 29.140 205.905 29.400 205.995 ;
        RECT 30.580 204.865 30.720 206.390 ;
        RECT 31.040 204.865 31.180 207.945 ;
        RECT 31.500 205.885 31.640 216.445 ;
        RECT 31.960 216.085 32.100 216.445 ;
        RECT 31.900 215.765 32.160 216.085 ;
        RECT 37.870 215.230 38.150 215.600 ;
        RECT 36.040 214.405 36.300 214.725 ;
        RECT 32.710 212.170 34.250 212.540 ;
        RECT 33.280 211.685 33.540 212.005 ;
        RECT 32.360 210.665 32.620 210.985 ;
        RECT 31.900 210.325 32.160 210.645 ;
        RECT 31.440 205.565 31.700 205.885 ;
        RECT 30.520 204.545 30.780 204.865 ;
        RECT 30.980 204.545 31.240 204.865 ;
        RECT 29.410 204.010 30.950 204.380 ;
        RECT 31.500 203.505 31.640 205.565 ;
        RECT 31.960 205.285 32.100 210.325 ;
        RECT 32.420 207.585 32.560 210.665 ;
        RECT 33.340 208.945 33.480 211.685 ;
        RECT 36.100 211.665 36.240 214.405 ;
        RECT 37.420 214.065 37.680 214.385 ;
        RECT 36.500 213.725 36.760 214.045 ;
        RECT 36.040 211.345 36.300 211.665 ;
        RECT 35.120 211.235 35.380 211.325 ;
        RECT 35.120 211.095 35.780 211.235 ;
        RECT 35.120 211.005 35.380 211.095 ;
        RECT 35.640 209.285 35.780 211.095 ;
        RECT 36.040 210.665 36.300 210.985 ;
        RECT 35.120 208.965 35.380 209.285 ;
        RECT 35.580 208.965 35.840 209.285 ;
        RECT 33.280 208.625 33.540 208.945 ;
        RECT 35.180 208.265 35.320 208.965 ;
        RECT 34.660 207.945 34.920 208.265 ;
        RECT 35.120 207.945 35.380 208.265 ;
        RECT 35.580 207.945 35.840 208.265 ;
        RECT 32.360 207.265 32.620 207.585 ;
        RECT 32.710 206.730 34.250 207.100 ;
        RECT 32.360 205.795 32.620 205.885 ;
        RECT 32.360 205.655 33.020 205.795 ;
        RECT 32.360 205.565 32.620 205.655 ;
        RECT 31.960 205.145 32.560 205.285 ;
        RECT 31.900 204.545 32.160 204.865 ;
        RECT 31.440 203.185 31.700 203.505 ;
        RECT 30.060 202.735 30.320 202.825 ;
        RECT 28.740 202.595 30.320 202.735 ;
        RECT 30.060 202.505 30.320 202.595 ;
        RECT 28.680 200.805 28.940 201.125 ;
        RECT 28.220 199.785 28.480 200.105 ;
        RECT 28.280 198.405 28.420 199.785 ;
        RECT 28.220 198.085 28.480 198.405 ;
        RECT 28.740 197.385 28.880 200.805 ;
        RECT 30.120 200.445 30.260 202.505 ;
        RECT 31.500 200.445 31.640 203.185 ;
        RECT 30.060 200.125 30.320 200.445 ;
        RECT 30.980 200.125 31.240 200.445 ;
        RECT 31.440 200.125 31.700 200.445 ;
        RECT 31.040 199.335 31.180 200.125 ;
        RECT 31.040 199.195 31.640 199.335 ;
        RECT 29.410 198.570 30.950 198.940 ;
        RECT 30.520 198.085 30.780 198.405 ;
        RECT 28.680 197.065 28.940 197.385 ;
        RECT 29.590 196.870 29.870 197.240 ;
        RECT 30.060 197.065 30.320 197.385 ;
        RECT 28.220 196.385 28.480 196.705 ;
        RECT 27.760 193.665 28.020 193.985 ;
        RECT 27.300 192.645 27.560 192.965 ;
        RECT 28.280 191.855 28.420 196.385 ;
        RECT 28.680 195.025 28.940 195.345 ;
        RECT 28.740 192.875 28.880 195.025 ;
        RECT 29.660 195.005 29.800 196.870 ;
        RECT 30.120 195.345 30.260 197.065 ;
        RECT 30.060 195.025 30.320 195.345 ;
        RECT 29.600 194.685 29.860 195.005 ;
        RECT 30.580 194.915 30.720 198.085 ;
        RECT 31.500 196.705 31.640 199.195 ;
        RECT 31.440 196.385 31.700 196.705 ;
        RECT 30.980 195.595 31.240 195.685 ;
        RECT 31.500 195.595 31.640 196.385 ;
        RECT 30.980 195.455 31.640 195.595 ;
        RECT 30.980 195.365 31.240 195.455 ;
        RECT 30.980 194.915 31.240 195.005 ;
        RECT 30.580 194.775 31.640 194.915 ;
        RECT 30.980 194.685 31.240 194.775 ;
        RECT 29.660 194.520 29.800 194.685 ;
        RECT 29.590 194.150 29.870 194.520 ;
        RECT 29.410 193.130 30.950 193.500 ;
        RECT 28.740 192.735 29.340 192.875 ;
        RECT 29.200 191.945 29.340 192.735 ;
        RECT 31.500 191.945 31.640 194.775 ;
        RECT 31.960 191.945 32.100 204.545 ;
        RECT 32.420 201.035 32.560 205.145 ;
        RECT 32.880 204.720 33.020 205.655 ;
        RECT 34.200 205.565 34.460 205.885 ;
        RECT 32.810 204.350 33.090 204.720 ;
        RECT 34.260 203.845 34.400 205.565 ;
        RECT 34.720 205.285 34.860 207.945 ;
        RECT 35.640 205.885 35.780 207.945 ;
        RECT 35.580 205.565 35.840 205.885 ;
        RECT 34.720 205.145 35.320 205.285 ;
        RECT 34.660 204.545 34.920 204.865 ;
        RECT 34.200 203.525 34.460 203.845 ;
        RECT 32.820 202.505 33.080 202.825 ;
        RECT 32.880 202.145 33.020 202.505 ;
        RECT 32.820 201.825 33.080 202.145 ;
        RECT 32.710 201.290 34.250 201.660 ;
        RECT 32.420 200.895 33.020 201.035 ;
        RECT 32.350 198.230 32.630 198.600 ;
        RECT 32.420 197.725 32.560 198.230 ;
        RECT 32.880 198.065 33.020 200.895 ;
        RECT 34.720 200.785 34.860 204.545 ;
        RECT 35.180 203.755 35.320 205.145 ;
        RECT 35.180 203.615 35.780 203.755 ;
        RECT 35.120 202.845 35.380 203.165 ;
        RECT 33.280 200.465 33.540 200.785 ;
        RECT 32.820 197.745 33.080 198.065 ;
        RECT 32.360 197.405 32.620 197.725 ;
        RECT 33.340 197.385 33.480 200.465 ;
        RECT 33.730 200.270 34.010 200.640 ;
        RECT 34.660 200.465 34.920 200.785 ;
        RECT 33.280 197.065 33.540 197.385 ;
        RECT 33.800 197.240 33.940 200.270 ;
        RECT 34.200 200.125 34.460 200.445 ;
        RECT 34.260 199.280 34.400 200.125 ;
        RECT 34.190 198.910 34.470 199.280 ;
        RECT 35.180 198.405 35.320 202.845 ;
        RECT 35.640 201.320 35.780 203.615 ;
        RECT 35.570 200.950 35.850 201.320 ;
        RECT 35.580 200.125 35.840 200.445 ;
        RECT 35.120 198.085 35.380 198.405 ;
        RECT 34.660 197.745 34.920 198.065 ;
        RECT 33.730 196.870 34.010 197.240 ;
        RECT 32.360 196.385 32.620 196.705 ;
        RECT 32.420 192.285 32.560 196.385 ;
        RECT 32.710 195.850 34.250 196.220 ;
        RECT 34.720 195.345 34.860 197.745 ;
        RECT 35.110 197.550 35.390 197.920 ;
        RECT 34.660 195.025 34.920 195.345 ;
        RECT 33.740 194.915 34.000 195.005 ;
        RECT 35.180 194.915 35.320 197.550 ;
        RECT 35.640 197.385 35.780 200.125 ;
        RECT 35.580 197.240 35.840 197.385 ;
        RECT 35.570 196.870 35.850 197.240 ;
        RECT 36.100 195.685 36.240 210.665 ;
        RECT 36.560 203.845 36.700 213.725 ;
        RECT 37.480 213.365 37.620 214.065 ;
        RECT 37.420 213.045 37.680 213.365 ;
        RECT 36.960 212.705 37.220 213.025 ;
        RECT 37.020 212.005 37.160 212.705 ;
        RECT 36.960 211.685 37.220 212.005 ;
        RECT 37.020 210.840 37.160 211.685 ;
        RECT 37.410 211.150 37.690 211.520 ;
        RECT 37.940 211.325 38.080 215.230 ;
        RECT 38.800 213.385 39.060 213.705 ;
        RECT 37.480 210.985 37.620 211.150 ;
        RECT 37.880 211.005 38.140 211.325 ;
        RECT 36.950 210.470 37.230 210.840 ;
        RECT 37.420 210.665 37.680 210.985 ;
        RECT 37.420 208.965 37.680 209.285 ;
        RECT 37.480 208.265 37.620 208.965 ;
        RECT 37.940 208.945 38.080 211.005 ;
        RECT 38.860 209.285 39.000 213.385 ;
        RECT 39.320 210.305 39.460 216.785 ;
        RECT 39.720 216.105 39.980 216.425 ;
        RECT 39.780 213.025 39.920 216.105 ;
        RECT 39.720 212.705 39.980 213.025 ;
        RECT 39.780 210.645 39.920 212.705 ;
        RECT 40.180 210.665 40.440 210.985 ;
        RECT 39.720 210.325 39.980 210.645 ;
        RECT 39.260 209.985 39.520 210.305 ;
        RECT 38.800 208.965 39.060 209.285 ;
        RECT 37.880 208.625 38.140 208.945 ;
        RECT 36.960 207.945 37.220 208.265 ;
        RECT 37.420 207.945 37.680 208.265 ;
        RECT 38.340 207.945 38.600 208.265 ;
        RECT 37.020 206.565 37.160 207.945 ;
        RECT 37.480 207.585 37.620 207.945 ;
        RECT 37.420 207.265 37.680 207.585 ;
        RECT 36.960 206.245 37.220 206.565 ;
        RECT 37.880 205.905 38.140 206.225 ;
        RECT 37.940 205.545 38.080 205.905 ;
        RECT 38.400 205.885 38.540 207.945 ;
        RECT 39.320 207.925 39.460 209.985 ;
        RECT 40.240 208.005 40.380 210.665 ;
        RECT 39.260 207.605 39.520 207.925 ;
        RECT 39.780 207.865 40.380 208.005 ;
        RECT 39.780 205.885 39.920 207.865 ;
        RECT 40.180 207.265 40.440 207.585 ;
        RECT 40.240 205.885 40.380 207.265 ;
        RECT 38.340 205.565 38.600 205.885 ;
        RECT 39.720 205.565 39.980 205.885 ;
        RECT 40.180 205.565 40.440 205.885 ;
        RECT 37.880 205.225 38.140 205.545 ;
        RECT 36.960 204.545 37.220 204.865 ;
        RECT 37.020 203.845 37.160 204.545 ;
        RECT 36.500 203.525 36.760 203.845 ;
        RECT 36.960 203.525 37.220 203.845 ;
        RECT 37.420 203.245 37.680 203.505 ;
        RECT 37.020 203.185 37.680 203.245 ;
        RECT 37.020 203.105 37.620 203.185 ;
        RECT 37.020 201.125 37.160 203.105 ;
        RECT 36.960 200.805 37.220 201.125 ;
        RECT 36.500 200.125 36.760 200.445 ;
        RECT 36.960 200.125 37.220 200.445 ;
        RECT 37.420 200.125 37.680 200.445 ;
        RECT 36.560 199.425 36.700 200.125 ;
        RECT 36.500 199.105 36.760 199.425 ;
        RECT 37.020 198.405 37.160 200.125 ;
        RECT 36.500 198.085 36.760 198.405 ;
        RECT 36.960 198.085 37.220 198.405 ;
        RECT 36.040 195.365 36.300 195.685 ;
        RECT 35.580 194.915 35.840 195.005 ;
        RECT 33.740 194.775 34.400 194.915 ;
        RECT 33.740 194.685 34.000 194.775 ;
        RECT 34.260 194.575 34.400 194.775 ;
        RECT 35.180 194.775 35.840 194.915 ;
        RECT 35.180 194.575 35.320 194.775 ;
        RECT 35.580 194.685 35.840 194.775 ;
        RECT 32.810 194.150 33.090 194.520 ;
        RECT 34.260 194.435 35.320 194.575 ;
        RECT 32.360 191.965 32.620 192.285 ;
        RECT 32.880 191.945 33.020 194.150 ;
        RECT 33.280 193.840 33.540 193.985 ;
        RECT 33.270 193.470 33.550 193.840 ;
        RECT 33.340 192.285 33.480 193.470 ;
        RECT 33.280 191.965 33.540 192.285 ;
        RECT 28.680 191.855 28.940 191.945 ;
        RECT 28.280 191.715 28.940 191.855 ;
        RECT 28.680 191.625 28.940 191.715 ;
        RECT 29.140 191.625 29.400 191.945 ;
        RECT 31.440 191.625 31.700 191.945 ;
        RECT 31.900 191.625 32.160 191.945 ;
        RECT 32.820 191.625 33.080 191.945 ;
        RECT 33.740 191.800 34.000 191.945 ;
        RECT 23.160 191.285 23.420 191.605 ;
        RECT 26.840 191.285 27.100 191.605 ;
        RECT 20.400 188.905 20.660 189.225 ;
        RECT 19.480 188.555 19.740 188.875 ;
        RECT 23.220 187.715 23.360 191.285 ;
        RECT 31.500 191.265 31.640 191.625 ;
        RECT 33.730 191.430 34.010 191.800 ;
        RECT 34.660 191.285 34.920 191.605 ;
        RECT 27.760 190.945 28.020 191.265 ;
        RECT 28.220 190.945 28.480 191.265 ;
        RECT 31.440 190.945 31.700 191.265 ;
        RECT 27.820 188.110 27.960 190.945 ;
        RECT 28.280 189.760 28.420 190.945 ;
        RECT 32.710 190.410 34.250 190.780 ;
        RECT 28.210 189.390 28.490 189.760 ;
        RECT 34.720 188.185 34.860 191.285 ;
        RECT 36.560 189.565 36.700 198.085 ;
        RECT 36.950 196.190 37.230 196.560 ;
        RECT 37.020 195.005 37.160 196.190 ;
        RECT 36.960 194.685 37.220 195.005 ;
        RECT 37.480 192.965 37.620 200.125 ;
        RECT 37.940 195.345 38.080 205.225 ;
        RECT 39.260 202.505 39.520 202.825 ;
        RECT 38.340 201.825 38.600 202.145 ;
        RECT 38.400 197.725 38.540 201.825 ;
        RECT 39.320 198.405 39.460 202.505 ;
        RECT 40.180 202.165 40.440 202.485 ;
        RECT 40.240 201.125 40.380 202.165 ;
        RECT 40.180 200.805 40.440 201.125 ;
        RECT 40.170 198.910 40.450 199.280 ;
        RECT 39.260 198.315 39.520 198.405 ;
        RECT 38.860 198.175 39.520 198.315 ;
        RECT 38.340 197.405 38.600 197.725 ;
        RECT 38.400 195.880 38.540 197.405 ;
        RECT 38.330 195.510 38.610 195.880 ;
        RECT 38.860 195.685 39.000 198.175 ;
        RECT 39.260 198.085 39.520 198.175 ;
        RECT 40.240 197.385 40.380 198.910 ;
        RECT 40.700 198.405 40.840 217.270 ;
        RECT 41.560 216.445 41.820 216.765 ;
        RECT 41.100 213.385 41.360 213.705 ;
        RECT 41.160 212.200 41.300 213.385 ;
        RECT 41.090 211.830 41.370 212.200 ;
        RECT 41.620 210.160 41.760 216.445 ;
        RECT 43.460 216.425 43.600 218.485 ;
        RECT 43.400 216.105 43.660 216.425 ;
        RECT 43.460 215.745 43.600 216.105 ;
        RECT 43.400 215.425 43.660 215.745 ;
        RECT 44.320 215.425 44.580 215.745 ;
        RECT 44.380 214.725 44.520 215.425 ;
        RECT 44.320 214.405 44.580 214.725 ;
        RECT 45.240 214.635 45.500 214.725 ;
        RECT 44.840 214.495 45.500 214.635 ;
        RECT 42.020 210.665 42.280 210.985 ;
        RECT 41.550 209.790 41.830 210.160 ;
        RECT 41.620 207.585 41.760 209.790 ;
        RECT 42.080 208.605 42.220 210.665 ;
        RECT 44.840 208.945 44.980 214.495 ;
        RECT 45.240 214.405 45.500 214.495 ;
        RECT 42.940 208.625 43.200 208.945 ;
        RECT 44.780 208.625 45.040 208.945 ;
        RECT 42.020 208.285 42.280 208.605 ;
        RECT 41.560 207.265 41.820 207.585 ;
        RECT 43.000 201.035 43.140 208.625 ;
        RECT 44.320 207.945 44.580 208.265 ;
        RECT 45.240 207.945 45.500 208.265 ;
        RECT 43.860 205.225 44.120 205.545 ;
        RECT 43.920 202.825 44.060 205.225 ;
        RECT 43.860 202.505 44.120 202.825 ;
        RECT 43.860 201.825 44.120 202.145 ;
        RECT 41.160 200.895 43.140 201.035 ;
        RECT 41.160 200.445 41.300 200.895 ;
        RECT 41.100 200.125 41.360 200.445 ;
        RECT 41.560 200.125 41.820 200.445 ;
        RECT 42.480 200.125 42.740 200.445 ;
        RECT 41.620 199.425 41.760 200.125 ;
        RECT 42.540 199.765 42.680 200.125 ;
        RECT 42.480 199.445 42.740 199.765 ;
        RECT 41.560 199.105 41.820 199.425 ;
        RECT 40.640 198.085 40.900 198.405 ;
        RECT 41.100 197.635 41.360 197.725 ;
        RECT 41.620 197.635 41.760 199.105 ;
        RECT 41.100 197.495 41.760 197.635 ;
        RECT 41.100 197.405 41.360 197.495 ;
        RECT 40.180 197.065 40.440 197.385 ;
        RECT 39.260 196.725 39.520 197.045 ;
        RECT 38.800 195.365 39.060 195.685 ;
        RECT 37.880 195.025 38.140 195.345 ;
        RECT 37.420 192.645 37.680 192.965 ;
        RECT 37.940 192.285 38.080 195.025 ;
        RECT 39.320 194.325 39.460 196.725 ;
        RECT 40.630 195.510 40.910 195.880 ;
        RECT 40.700 195.005 40.840 195.510 ;
        RECT 41.160 195.005 41.300 197.405 ;
        RECT 43.000 197.385 43.140 200.895 ;
        RECT 43.920 199.765 44.060 201.825 ;
        RECT 43.400 199.445 43.660 199.765 ;
        RECT 43.860 199.445 44.120 199.765 ;
        RECT 43.460 197.725 43.600 199.445 ;
        RECT 44.380 199.280 44.520 207.945 ;
        RECT 45.300 207.440 45.440 207.945 ;
        RECT 45.230 207.070 45.510 207.440 ;
        RECT 45.760 204.720 45.900 219.165 ;
        RECT 49.380 218.485 49.640 218.805 ;
        RECT 46.160 216.785 46.420 217.105 ;
        RECT 46.220 216.280 46.360 216.785 ;
        RECT 46.150 215.910 46.430 216.280 ;
        RECT 46.620 216.105 46.880 216.425 ;
        RECT 47.080 216.105 47.340 216.425 ;
        RECT 46.680 212.005 46.820 216.105 ;
        RECT 46.620 211.685 46.880 212.005 ;
        RECT 47.140 209.285 47.280 216.105 ;
        RECT 48.920 211.685 49.180 212.005 ;
        RECT 48.980 211.325 49.120 211.685 ;
        RECT 48.920 211.005 49.180 211.325 ;
        RECT 47.540 209.985 47.800 210.305 ;
        RECT 47.080 208.965 47.340 209.285 ;
        RECT 46.620 207.945 46.880 208.265 ;
        RECT 46.150 205.710 46.430 206.080 ;
        RECT 46.680 205.885 46.820 207.945 ;
        RECT 47.600 207.585 47.740 209.985 ;
        RECT 49.440 208.265 49.580 218.485 ;
        RECT 50.750 218.265 51.030 219.340 ;
        RECT 59.960 218.825 60.220 219.145 ;
        RECT 50.820 217.445 50.960 218.265 ;
        RECT 50.760 217.125 51.020 217.445 ;
        RECT 53.520 216.785 53.780 217.105 ;
        RECT 53.580 214.725 53.720 216.785 ;
        RECT 55.350 215.910 55.630 216.280 ;
        RECT 57.200 216.105 57.460 216.425 ;
        RECT 53.520 214.405 53.780 214.725 ;
        RECT 54.900 214.405 55.160 214.725 ;
        RECT 49.840 212.705 50.100 213.025 ;
        RECT 49.900 211.325 50.040 212.705 ;
        RECT 51.680 211.345 51.940 211.665 ;
        RECT 49.840 211.005 50.100 211.325 ;
        RECT 50.760 211.005 51.020 211.325 ;
        RECT 48.000 207.945 48.260 208.265 ;
        RECT 49.380 207.945 49.640 208.265 ;
        RECT 47.540 207.265 47.800 207.585 ;
        RECT 45.690 204.350 45.970 204.720 ;
        RECT 45.240 203.525 45.500 203.845 ;
        RECT 45.300 202.825 45.440 203.525 ;
        RECT 45.240 202.505 45.500 202.825 ;
        RECT 44.780 201.825 45.040 202.145 ;
        RECT 44.310 198.910 44.590 199.280 ;
        RECT 44.840 198.600 44.980 201.825 ;
        RECT 45.760 201.125 45.900 204.350 ;
        RECT 45.700 200.805 45.960 201.125 ;
        RECT 45.240 200.465 45.500 200.785 ;
        RECT 45.300 199.960 45.440 200.465 ;
        RECT 45.700 200.125 45.960 200.445 ;
        RECT 45.230 199.590 45.510 199.960 ;
        RECT 44.770 198.230 45.050 198.600 ;
        RECT 43.400 197.405 43.660 197.725 ;
        RECT 42.940 197.065 43.200 197.385 ;
        RECT 43.000 196.705 43.140 197.065 ;
        RECT 42.940 196.385 43.200 196.705 ;
        RECT 43.460 195.685 43.600 197.405 ;
        RECT 45.760 197.385 45.900 200.125 ;
        RECT 46.220 197.920 46.360 205.710 ;
        RECT 46.620 205.565 46.880 205.885 ;
        RECT 47.070 205.710 47.350 206.080 ;
        RECT 47.140 205.545 47.280 205.710 ;
        RECT 47.080 205.225 47.340 205.545 ;
        RECT 46.620 202.735 46.880 202.825 ;
        RECT 47.600 202.735 47.740 207.265 ;
        RECT 48.060 205.885 48.200 207.945 ;
        RECT 48.920 205.905 49.180 206.225 ;
        RECT 48.000 205.565 48.260 205.885 ;
        RECT 48.060 205.205 48.200 205.565 ;
        RECT 48.000 204.885 48.260 205.205 ;
        RECT 48.060 202.825 48.200 204.885 ;
        RECT 48.980 202.825 49.120 205.905 ;
        RECT 49.440 205.885 49.580 207.945 ;
        RECT 49.900 206.565 50.040 211.005 ;
        RECT 50.290 208.430 50.570 208.800 ;
        RECT 50.360 208.265 50.500 208.430 ;
        RECT 50.300 207.945 50.560 208.265 ;
        RECT 50.290 207.070 50.570 207.440 ;
        RECT 49.840 206.245 50.100 206.565 ;
        RECT 49.380 205.565 49.640 205.885 ;
        RECT 49.830 205.710 50.110 206.080 ;
        RECT 49.840 205.565 50.100 205.710 ;
        RECT 49.380 204.545 49.640 204.865 ;
        RECT 46.620 202.595 47.740 202.735 ;
        RECT 46.620 202.505 46.880 202.595 ;
        RECT 48.000 202.505 48.260 202.825 ;
        RECT 48.920 202.505 49.180 202.825 ;
        RECT 46.150 197.550 46.430 197.920 ;
        RECT 45.700 197.065 45.960 197.385 ;
        RECT 46.680 195.880 46.820 202.505 ;
        RECT 48.060 202.000 48.200 202.505 ;
        RECT 49.440 202.485 49.580 204.545 ;
        RECT 48.460 202.165 48.720 202.485 ;
        RECT 49.380 202.165 49.640 202.485 ;
        RECT 47.990 201.630 48.270 202.000 ;
        RECT 48.520 201.125 48.660 202.165 ;
        RECT 48.460 201.035 48.720 201.125 ;
        RECT 48.060 200.895 48.720 201.035 ;
        RECT 48.060 200.525 48.200 200.895 ;
        RECT 48.460 200.805 48.720 200.895 ;
        RECT 47.140 200.385 48.200 200.525 ;
        RECT 47.140 197.045 47.280 200.385 ;
        RECT 48.460 200.355 48.720 200.445 ;
        RECT 49.440 200.355 49.580 202.165 ;
        RECT 48.460 200.215 49.580 200.355 ;
        RECT 48.460 200.125 48.720 200.215 ;
        RECT 47.540 199.785 47.800 200.105 ;
        RECT 47.080 196.725 47.340 197.045 ;
        RECT 43.400 195.365 43.660 195.685 ;
        RECT 46.610 195.510 46.890 195.880 ;
        RECT 41.560 195.025 41.820 195.345 ;
        RECT 40.640 194.685 40.900 195.005 ;
        RECT 41.100 194.685 41.360 195.005 ;
        RECT 39.260 194.005 39.520 194.325 ;
        RECT 40.640 193.665 40.900 193.985 ;
        RECT 38.340 192.645 38.600 192.965 ;
        RECT 37.880 191.965 38.140 192.285 ;
        RECT 38.400 190.185 38.540 192.645 ;
        RECT 40.700 192.625 40.840 193.665 ;
        RECT 41.620 192.965 41.760 195.025 ;
        RECT 47.600 195.005 47.740 199.785 ;
        RECT 48.000 199.105 48.260 199.425 ;
        RECT 47.540 194.685 47.800 195.005 ;
        RECT 48.060 194.665 48.200 199.105 ;
        RECT 48.520 195.685 48.660 200.125 ;
        RECT 48.920 198.085 49.180 198.405 ;
        RECT 48.980 197.725 49.120 198.085 ;
        RECT 48.920 197.405 49.180 197.725 ;
        RECT 48.980 197.240 49.120 197.405 ;
        RECT 48.910 196.870 49.190 197.240 ;
        RECT 49.380 196.725 49.640 197.045 ;
        RECT 48.920 196.385 49.180 196.705 ;
        RECT 48.460 195.365 48.720 195.685 ;
        RECT 43.400 194.345 43.660 194.665 ;
        RECT 48.000 194.345 48.260 194.665 ;
        RECT 41.560 192.645 41.820 192.965 ;
        RECT 40.640 192.305 40.900 192.625 ;
        RECT 43.460 192.285 43.600 194.345 ;
        RECT 47.080 193.665 47.340 193.985 ;
        RECT 43.400 191.965 43.660 192.285 ;
        RECT 38.800 191.625 39.060 191.945 ;
        RECT 41.560 191.625 41.820 191.945 ;
        RECT 38.860 190.245 39.000 191.625 ;
        RECT 37.020 190.045 38.540 190.185 ;
        RECT 37.020 189.660 37.160 190.045 ;
        RECT 38.800 189.925 39.060 190.245 ;
        RECT 41.620 189.660 41.760 191.625 ;
        RECT 46.160 190.945 46.420 191.265 ;
        RECT 36.500 189.245 36.760 189.565 ;
        RECT 37.020 189.520 41.760 189.660 ;
        RECT 32.360 188.110 32.620 188.185 ;
        RECT 27.820 187.970 32.620 188.110 ;
        RECT 27.820 187.715 27.960 187.970 ;
        RECT 32.360 187.865 32.620 187.970 ;
        RECT 34.660 187.865 34.920 188.185 ;
        RECT 32.420 187.715 32.560 187.865 ;
        RECT 37.020 187.715 37.160 189.520 ;
        RECT 41.620 187.715 41.760 189.520 ;
        RECT 46.220 188.960 46.360 190.945 ;
        RECT 47.140 189.905 47.280 193.665 ;
        RECT 48.520 191.945 48.660 195.365 ;
        RECT 48.460 191.625 48.720 191.945 ;
        RECT 47.540 190.945 47.800 191.265 ;
        RECT 47.600 189.905 47.740 190.945 ;
        RECT 47.080 189.585 47.340 189.905 ;
        RECT 47.540 189.585 47.800 189.905 ;
        RECT 48.980 189.760 49.120 196.385 ;
        RECT 49.440 190.440 49.580 196.725 ;
        RECT 49.900 192.625 50.040 205.565 ;
        RECT 50.360 203.415 50.500 207.070 ;
        RECT 50.820 204.865 50.960 211.005 ;
        RECT 51.220 209.985 51.480 210.305 ;
        RECT 50.760 204.545 51.020 204.865 ;
        RECT 50.760 203.415 51.020 203.505 ;
        RECT 50.360 203.275 51.020 203.415 ;
        RECT 50.760 203.185 51.020 203.275 ;
        RECT 50.820 202.825 50.960 203.185 ;
        RECT 50.760 202.505 51.020 202.825 ;
        RECT 50.290 200.950 50.570 201.320 ;
        RECT 50.360 199.765 50.500 200.950 ;
        RECT 50.300 199.445 50.560 199.765 ;
        RECT 50.360 199.280 50.500 199.445 ;
        RECT 50.290 198.910 50.570 199.280 ;
        RECT 50.290 198.230 50.570 198.600 ;
        RECT 50.360 195.345 50.500 198.230 ;
        RECT 50.760 197.405 51.020 197.725 ;
        RECT 50.300 195.025 50.560 195.345 ;
        RECT 49.840 192.305 50.100 192.625 ;
        RECT 49.900 191.945 50.040 192.305 ;
        RECT 49.840 191.625 50.100 191.945 ;
        RECT 49.370 190.070 49.650 190.440 ;
        RECT 48.910 189.390 49.190 189.760 ;
        RECT 50.820 188.960 50.960 197.405 ;
        RECT 46.220 188.820 50.960 188.960 ;
        RECT 46.220 187.715 46.360 188.820 ;
        RECT 50.820 187.715 50.960 188.820 ;
        RECT 51.280 188.545 51.420 209.985 ;
        RECT 51.740 207.585 51.880 211.345 ;
        RECT 52.140 211.005 52.400 211.325 ;
        RECT 52.200 209.285 52.340 211.005 ;
        RECT 53.060 209.985 53.320 210.305 ;
        RECT 52.140 208.965 52.400 209.285 ;
        RECT 53.120 208.605 53.260 209.985 ;
        RECT 53.580 209.285 53.720 214.405 ;
        RECT 54.960 212.005 55.100 214.405 ;
        RECT 54.900 211.685 55.160 212.005 ;
        RECT 54.890 211.150 55.170 211.520 ;
        RECT 55.420 211.325 55.560 215.910 ;
        RECT 56.740 214.405 57.000 214.725 ;
        RECT 56.800 213.365 56.940 214.405 ;
        RECT 56.740 213.045 57.000 213.365 ;
        RECT 56.740 211.685 57.000 212.005 ;
        RECT 54.960 210.985 55.100 211.150 ;
        RECT 55.360 211.005 55.620 211.325 ;
        RECT 54.900 210.665 55.160 210.985 ;
        RECT 55.820 210.665 56.080 210.985 ;
        RECT 55.360 210.325 55.620 210.645 ;
        RECT 53.520 208.965 53.780 209.285 ;
        RECT 54.890 209.110 55.170 209.480 ;
        RECT 53.060 208.285 53.320 208.605 ;
        RECT 53.050 207.750 53.330 208.120 ;
        RECT 51.680 207.265 51.940 207.585 ;
        RECT 51.740 205.205 51.880 207.265 ;
        RECT 51.680 204.885 51.940 205.205 ;
        RECT 51.680 199.785 51.940 200.105 ;
        RECT 52.600 199.960 52.860 200.105 ;
        RECT 51.740 198.405 51.880 199.785 ;
        RECT 52.590 199.590 52.870 199.960 ;
        RECT 51.680 198.085 51.940 198.405 ;
        RECT 53.120 197.385 53.260 207.750 ;
        RECT 53.520 205.565 53.780 205.885 ;
        RECT 53.970 205.710 54.250 206.080 ;
        RECT 53.980 205.565 54.240 205.710 ;
        RECT 54.440 205.565 54.700 205.885 ;
        RECT 53.580 200.785 53.720 205.565 ;
        RECT 53.980 204.545 54.240 204.865 ;
        RECT 53.520 200.465 53.780 200.785 ;
        RECT 51.680 197.065 51.940 197.385 ;
        RECT 51.740 195.685 51.880 197.065 ;
        RECT 52.140 196.725 52.400 197.045 ;
        RECT 52.590 196.870 52.870 197.240 ;
        RECT 53.060 197.065 53.320 197.385 ;
        RECT 52.200 195.685 52.340 196.725 ;
        RECT 51.680 195.365 51.940 195.685 ;
        RECT 52.140 195.365 52.400 195.685 ;
        RECT 52.140 194.685 52.400 195.005 ;
        RECT 52.200 191.945 52.340 194.685 ;
        RECT 52.660 194.665 52.800 196.870 ;
        RECT 53.060 196.385 53.320 196.705 ;
        RECT 52.600 194.345 52.860 194.665 ;
        RECT 51.670 191.430 51.950 191.800 ;
        RECT 52.140 191.625 52.400 191.945 ;
        RECT 52.660 191.605 52.800 194.345 ;
        RECT 53.120 192.625 53.260 196.385 ;
        RECT 53.580 195.005 53.720 200.465 ;
        RECT 53.520 194.685 53.780 195.005 ;
        RECT 53.580 193.985 53.720 194.685 ;
        RECT 53.520 193.665 53.780 193.985 ;
        RECT 53.060 192.305 53.320 192.625 ;
        RECT 51.740 191.265 51.880 191.430 ;
        RECT 52.600 191.285 52.860 191.605 ;
        RECT 51.680 190.945 51.940 191.265 ;
        RECT 54.040 188.885 54.180 204.545 ;
        RECT 54.500 203.505 54.640 205.565 ;
        RECT 54.440 203.185 54.700 203.505 ;
        RECT 54.500 199.280 54.640 203.185 ;
        RECT 54.430 198.910 54.710 199.280 ;
        RECT 54.960 198.405 55.100 209.110 ;
        RECT 55.420 208.265 55.560 210.325 ;
        RECT 55.880 209.285 56.020 210.665 ;
        RECT 56.270 209.790 56.550 210.160 ;
        RECT 56.340 209.285 56.480 209.790 ;
        RECT 55.820 208.965 56.080 209.285 ;
        RECT 56.280 208.965 56.540 209.285 ;
        RECT 56.800 208.265 56.940 211.685 ;
        RECT 57.260 211.665 57.400 216.105 ;
        RECT 58.120 215.425 58.380 215.745 ;
        RECT 57.200 211.345 57.460 211.665 ;
        RECT 55.360 207.945 55.620 208.265 ;
        RECT 56.740 207.945 57.000 208.265 ;
        RECT 57.260 206.080 57.400 211.345 ;
        RECT 57.660 210.665 57.920 210.985 ;
        RECT 57.720 206.565 57.860 210.665 ;
        RECT 58.180 206.565 58.320 215.425 ;
        RECT 59.040 208.625 59.300 208.945 ;
        RECT 57.660 206.245 57.920 206.565 ;
        RECT 58.120 206.245 58.380 206.565 ;
        RECT 55.810 205.710 56.090 206.080 ;
        RECT 56.280 205.795 56.540 205.885 ;
        RECT 55.880 203.505 56.020 205.710 ;
        RECT 56.280 205.655 56.940 205.795 ;
        RECT 57.190 205.710 57.470 206.080 ;
        RECT 58.580 205.905 58.840 206.225 ;
        RECT 56.280 205.565 56.540 205.655 ;
        RECT 56.800 205.455 56.940 205.655 ;
        RECT 57.200 205.455 57.460 205.545 ;
        RECT 56.800 205.315 57.460 205.455 ;
        RECT 55.820 203.185 56.080 203.505 ;
        RECT 55.360 200.125 55.620 200.445 ;
        RECT 54.900 198.085 55.160 198.405 ;
        RECT 55.420 196.705 55.560 200.125 ;
        RECT 55.880 198.485 56.020 203.185 ;
        RECT 56.280 202.505 56.540 202.825 ;
        RECT 56.800 202.735 56.940 205.315 ;
        RECT 57.200 205.225 57.460 205.315 ;
        RECT 58.120 204.885 58.380 205.205 ;
        RECT 58.180 204.040 58.320 204.885 ;
        RECT 58.110 203.670 58.390 204.040 ;
        RECT 58.180 202.825 58.320 203.670 ;
        RECT 58.640 202.825 58.780 205.905 ;
        RECT 59.100 202.825 59.240 208.625 ;
        RECT 59.500 207.265 59.760 207.585 ;
        RECT 59.560 205.205 59.700 207.265 ;
        RECT 59.500 204.885 59.760 205.205 ;
        RECT 57.200 202.735 57.460 202.825 ;
        RECT 56.800 202.595 57.460 202.735 ;
        RECT 57.200 202.505 57.460 202.595 ;
        RECT 58.120 202.505 58.380 202.825 ;
        RECT 58.580 202.505 58.840 202.825 ;
        RECT 59.040 202.505 59.300 202.825 ;
        RECT 56.340 199.425 56.480 202.505 ;
        RECT 57.260 202.145 57.400 202.505 ;
        RECT 57.200 201.825 57.460 202.145 ;
        RECT 56.730 200.950 57.010 201.320 ;
        RECT 56.800 200.445 56.940 200.950 ;
        RECT 56.740 200.125 57.000 200.445 ;
        RECT 56.730 199.590 57.010 199.960 ;
        RECT 56.740 199.445 57.000 199.590 ;
        RECT 56.280 199.105 56.540 199.425 ;
        RECT 55.880 198.345 56.940 198.485 ;
        RECT 56.280 197.405 56.540 197.725 ;
        RECT 55.360 196.385 55.620 196.705 ;
        RECT 54.890 195.510 55.170 195.880 ;
        RECT 54.900 195.365 55.160 195.510 ;
        RECT 54.960 194.325 55.100 195.365 ;
        RECT 55.420 195.005 55.560 196.385 ;
        RECT 55.820 195.365 56.080 195.685 ;
        RECT 55.360 194.685 55.620 195.005 ;
        RECT 54.900 194.005 55.160 194.325 ;
        RECT 55.880 193.985 56.020 195.365 ;
        RECT 56.340 195.345 56.480 197.405 ;
        RECT 56.280 195.025 56.540 195.345 ;
        RECT 55.820 193.665 56.080 193.985 ;
        RECT 55.820 192.875 56.080 192.965 ;
        RECT 56.340 192.875 56.480 195.025 ;
        RECT 55.820 192.735 56.480 192.875 ;
        RECT 55.820 192.645 56.080 192.735 ;
        RECT 55.820 191.625 56.080 191.945 ;
        RECT 54.440 191.120 54.700 191.265 ;
        RECT 54.430 190.750 54.710 191.120 ;
        RECT 55.360 190.945 55.620 191.265 ;
        RECT 53.980 188.565 54.240 188.885 ;
        RECT 51.220 188.225 51.480 188.545 ;
        RECT 55.420 187.715 55.560 190.945 ;
        RECT 55.880 188.205 56.020 191.625 ;
        RECT 56.280 191.515 56.540 191.605 ;
        RECT 56.800 191.515 56.940 198.345 ;
        RECT 57.260 195.765 57.400 201.825 ;
        RECT 57.660 200.525 57.920 200.785 ;
        RECT 58.640 200.525 58.780 202.505 ;
        RECT 57.660 200.465 58.780 200.525 ;
        RECT 57.720 200.385 58.780 200.465 ;
        RECT 58.120 199.445 58.380 199.765 ;
        RECT 57.650 198.230 57.930 198.600 ;
        RECT 58.180 198.405 58.320 199.445 ;
        RECT 58.640 198.405 58.780 200.385 ;
        RECT 57.720 196.705 57.860 198.230 ;
        RECT 58.120 198.085 58.380 198.405 ;
        RECT 58.580 198.085 58.840 198.405 ;
        RECT 59.100 197.805 59.240 202.505 ;
        RECT 60.020 201.035 60.160 218.825 ;
        RECT 62.710 218.265 62.990 220.625 ;
        RECT 74.650 220.025 74.950 220.425 ;
        RECT 65.020 218.485 65.280 218.805 ;
        RECT 62.780 217.445 62.920 218.265 ;
        RECT 62.720 217.125 62.980 217.445 ;
        RECT 64.560 216.785 64.820 217.105 ;
        RECT 62.720 216.445 62.980 216.765 ;
        RECT 62.260 216.105 62.520 216.425 ;
        RECT 60.880 215.425 61.140 215.745 ;
        RECT 60.940 214.725 61.080 215.425 ;
        RECT 62.320 214.725 62.460 216.105 ;
        RECT 62.780 214.725 62.920 216.445 ;
        RECT 60.880 214.405 61.140 214.725 ;
        RECT 62.260 214.405 62.520 214.725 ;
        RECT 62.720 214.405 62.980 214.725 ;
        RECT 64.100 214.405 64.360 214.725 ;
        RECT 60.940 213.705 61.080 214.405 ;
        RECT 60.880 213.385 61.140 213.705 ;
        RECT 63.640 213.385 63.900 213.705 ;
        RECT 61.340 212.705 61.600 213.025 ;
        RECT 61.400 212.005 61.540 212.705 ;
        RECT 62.250 212.510 62.530 212.880 ;
        RECT 62.320 212.005 62.460 212.510 ;
        RECT 61.340 211.685 61.600 212.005 ;
        RECT 62.260 211.915 62.520 212.005 ;
        RECT 61.860 211.775 62.520 211.915 ;
        RECT 60.880 211.345 61.140 211.665 ;
        RECT 60.940 210.985 61.080 211.345 ;
        RECT 60.880 210.665 61.140 210.985 ;
        RECT 61.400 208.945 61.540 211.685 ;
        RECT 61.340 208.625 61.600 208.945 ;
        RECT 60.880 206.245 61.140 206.565 ;
        RECT 60.940 202.825 61.080 206.245 ;
        RECT 61.860 206.225 62.000 211.775 ;
        RECT 62.260 211.685 62.520 211.775 ;
        RECT 63.180 210.665 63.440 210.985 ;
        RECT 63.240 208.605 63.380 210.665 ;
        RECT 63.180 208.285 63.440 208.605 ;
        RECT 61.800 205.905 62.060 206.225 ;
        RECT 62.250 205.710 62.530 206.080 ;
        RECT 63.240 205.885 63.380 208.285 ;
        RECT 62.260 205.565 62.520 205.710 ;
        RECT 63.180 205.565 63.440 205.885 ;
        RECT 61.340 205.225 61.600 205.545 ;
        RECT 61.400 202.825 61.540 205.225 ;
        RECT 60.880 202.505 61.140 202.825 ;
        RECT 61.340 202.505 61.600 202.825 ;
        RECT 61.400 201.125 61.540 202.505 ;
        RECT 62.720 201.825 62.980 202.145 ;
        RECT 59.560 200.895 60.160 201.035 ;
        RECT 59.560 198.600 59.700 200.895 ;
        RECT 61.340 200.805 61.600 201.125 ;
        RECT 61.800 200.525 62.060 200.785 ;
        RECT 61.800 200.465 62.460 200.525 ;
        RECT 59.960 200.125 60.220 200.445 ;
        RECT 61.860 200.385 62.460 200.465 ;
        RECT 62.780 200.445 62.920 201.825 ;
        RECT 60.020 199.960 60.160 200.125 ;
        RECT 59.950 199.590 60.230 199.960 ;
        RECT 61.800 199.785 62.060 200.105 ;
        RECT 59.490 198.230 59.770 198.600 ;
        RECT 58.180 197.665 59.240 197.805 ;
        RECT 58.180 197.385 58.320 197.665 ;
        RECT 58.120 197.065 58.380 197.385 ;
        RECT 59.040 197.065 59.300 197.385 ;
        RECT 59.500 197.065 59.760 197.385 ;
        RECT 57.660 196.385 57.920 196.705 ;
        RECT 58.120 196.385 58.380 196.705 ;
        RECT 58.180 195.765 58.320 196.385 ;
        RECT 57.260 195.625 58.320 195.765 ;
        RECT 59.100 195.685 59.240 197.065 ;
        RECT 59.560 195.685 59.700 197.065 ;
        RECT 61.340 196.725 61.600 197.045 ;
        RECT 61.400 195.685 61.540 196.725 ;
        RECT 57.260 192.285 57.400 195.625 ;
        RECT 58.180 195.345 58.320 195.625 ;
        RECT 59.040 195.365 59.300 195.685 ;
        RECT 59.500 195.365 59.760 195.685 ;
        RECT 61.340 195.365 61.600 195.685 ;
        RECT 58.120 195.025 58.380 195.345 ;
        RECT 59.040 194.915 59.300 195.005 ;
        RECT 59.040 194.775 59.700 194.915 ;
        RECT 59.040 194.685 59.300 194.775 ;
        RECT 59.560 194.325 59.700 194.775 ;
        RECT 60.420 194.685 60.680 195.005 ;
        RECT 60.480 194.520 60.620 194.685 ;
        RECT 59.500 194.005 59.760 194.325 ;
        RECT 60.410 194.150 60.690 194.520 ;
        RECT 58.120 193.665 58.380 193.985 ;
        RECT 57.200 191.965 57.460 192.285 ;
        RECT 57.660 191.795 57.920 192.115 ;
        RECT 57.720 191.515 57.860 191.795 ;
        RECT 56.280 191.375 57.860 191.515 ;
        RECT 56.280 191.285 56.540 191.375 ;
        RECT 58.180 188.545 58.320 193.665 ;
        RECT 58.580 191.625 58.840 191.945 ;
        RECT 59.960 191.625 60.220 191.945 ;
        RECT 58.640 191.120 58.780 191.625 ;
        RECT 58.570 190.750 58.850 191.120 ;
        RECT 58.120 188.225 58.380 188.545 ;
        RECT 55.820 187.885 56.080 188.205 ;
        RECT 60.020 187.715 60.160 191.625 ;
        RECT 60.420 190.945 60.680 191.265 ;
        RECT 60.480 188.205 60.620 190.945 ;
        RECT 61.860 189.225 62.000 199.785 ;
        RECT 62.320 199.765 62.460 200.385 ;
        RECT 62.720 200.125 62.980 200.445 ;
        RECT 63.700 200.105 63.840 213.385 ;
        RECT 64.160 207.925 64.300 214.405 ;
        RECT 64.620 212.005 64.760 216.785 ;
        RECT 65.080 214.045 65.220 218.485 ;
        RECT 74.670 218.265 74.950 220.025 ;
        RECT 86.630 219.850 86.910 220.265 ;
        RECT 86.610 219.450 86.910 219.850 ;
        RECT 84.340 218.485 84.600 218.805 ;
        RECT 74.740 217.445 74.880 218.265 ;
        RECT 74.680 217.125 74.940 217.445 ;
        RECT 70.540 216.785 70.800 217.105 ;
        RECT 77.440 216.785 77.700 217.105 ;
        RECT 70.080 216.445 70.340 216.765 ;
        RECT 65.470 215.910 65.750 216.280 ;
        RECT 69.160 216.105 69.420 216.425 ;
        RECT 65.020 213.725 65.280 214.045 ;
        RECT 64.560 211.685 64.820 212.005 ;
        RECT 64.100 207.605 64.360 207.925 ;
        RECT 65.540 206.225 65.680 215.910 ;
        RECT 68.690 214.550 68.970 214.920 ;
        RECT 66.860 213.385 67.120 213.705 ;
        RECT 65.940 211.345 66.200 211.665 ;
        RECT 65.480 205.905 65.740 206.225 ;
        RECT 64.100 205.565 64.360 205.885 ;
        RECT 65.020 205.565 65.280 205.885 ;
        RECT 64.160 203.505 64.300 205.565 ;
        RECT 65.080 205.205 65.220 205.565 ;
        RECT 65.020 204.885 65.280 205.205 ;
        RECT 64.100 203.185 64.360 203.505 ;
        RECT 64.160 200.445 64.300 203.185 ;
        RECT 65.080 201.125 65.220 204.885 ;
        RECT 66.000 203.505 66.140 211.345 ;
        RECT 66.920 208.605 67.060 213.385 ;
        RECT 68.240 213.045 68.500 213.365 ;
        RECT 68.300 212.005 68.440 213.045 ;
        RECT 68.240 211.685 68.500 212.005 ;
        RECT 67.780 211.005 68.040 211.325 ;
        RECT 66.860 208.285 67.120 208.605 ;
        RECT 66.400 207.605 66.660 207.925 ;
        RECT 66.460 205.205 66.600 207.605 ;
        RECT 66.400 204.885 66.660 205.205 ;
        RECT 66.920 203.845 67.060 208.285 ;
        RECT 67.840 206.225 67.980 211.005 ;
        RECT 68.760 209.285 68.900 214.550 ;
        RECT 69.220 211.575 69.360 216.105 ;
        RECT 69.620 211.575 69.880 211.665 ;
        RECT 69.220 211.435 69.880 211.575 ;
        RECT 69.220 210.305 69.360 211.435 ;
        RECT 69.620 211.345 69.880 211.435 ;
        RECT 70.140 210.985 70.280 216.445 ;
        RECT 70.600 215.745 70.740 216.785 ;
        RECT 70.540 215.425 70.800 215.745 ;
        RECT 71.000 215.425 71.260 215.745 ;
        RECT 71.060 212.005 71.200 215.425 ;
        RECT 71.920 213.955 72.180 214.045 ;
        RECT 71.920 213.815 73.040 213.955 ;
        RECT 71.920 213.725 72.180 213.815 ;
        RECT 71.450 213.190 71.730 213.560 ;
        RECT 72.370 213.190 72.650 213.560 ;
        RECT 71.000 211.685 71.260 212.005 ;
        RECT 70.080 210.665 70.340 210.985 ;
        RECT 69.160 209.985 69.420 210.305 ;
        RECT 70.080 209.985 70.340 210.305 ;
        RECT 68.700 208.965 68.960 209.285 ;
        RECT 70.140 208.605 70.280 209.985 ;
        RECT 70.530 209.110 70.810 209.480 ;
        RECT 71.520 209.285 71.660 213.190 ;
        RECT 72.440 213.025 72.580 213.190 ;
        RECT 72.380 212.705 72.640 213.025 ;
        RECT 71.920 210.325 72.180 210.645 ;
        RECT 71.980 209.285 72.120 210.325 ;
        RECT 72.370 209.790 72.650 210.160 ;
        RECT 70.080 208.285 70.340 208.605 ;
        RECT 67.780 205.905 68.040 206.225 ;
        RECT 69.620 205.905 69.880 206.225 ;
        RECT 68.700 205.225 68.960 205.545 ;
        RECT 67.320 204.545 67.580 204.865 ;
        RECT 66.400 203.525 66.660 203.845 ;
        RECT 66.860 203.525 67.120 203.845 ;
        RECT 65.940 203.185 66.200 203.505 ;
        RECT 66.460 203.165 66.600 203.525 ;
        RECT 66.400 202.845 66.660 203.165 ;
        RECT 65.020 200.805 65.280 201.125 ;
        RECT 64.100 200.125 64.360 200.445 ;
        RECT 63.640 199.785 63.900 200.105 ;
        RECT 66.400 199.785 66.660 200.105 ;
        RECT 62.260 199.445 62.520 199.765 ;
        RECT 63.180 198.085 63.440 198.405 ;
        RECT 62.260 195.365 62.520 195.685 ;
        RECT 62.710 195.510 62.990 195.880 ;
        RECT 62.320 193.985 62.460 195.365 ;
        RECT 62.260 193.665 62.520 193.985 ;
        RECT 62.780 191.945 62.920 195.510 ;
        RECT 63.240 194.325 63.380 198.085 ;
        RECT 66.460 197.385 66.600 199.785 ;
        RECT 66.920 198.065 67.060 203.525 ;
        RECT 67.380 202.825 67.520 204.545 ;
        RECT 67.320 202.505 67.580 202.825 ;
        RECT 68.240 201.825 68.500 202.145 ;
        RECT 68.300 200.445 68.440 201.825 ;
        RECT 68.760 201.125 68.900 205.225 ;
        RECT 69.160 202.165 69.420 202.485 ;
        RECT 69.220 201.125 69.360 202.165 ;
        RECT 68.700 200.805 68.960 201.125 ;
        RECT 69.160 200.805 69.420 201.125 ;
        RECT 69.680 201.035 69.820 205.905 ;
        RECT 70.080 205.795 70.340 205.885 ;
        RECT 70.600 205.795 70.740 209.110 ;
        RECT 71.460 208.965 71.720 209.285 ;
        RECT 71.920 208.965 72.180 209.285 ;
        RECT 72.440 208.605 72.580 209.790 ;
        RECT 72.380 208.285 72.640 208.605 ;
        RECT 70.080 205.655 70.740 205.795 ;
        RECT 70.080 205.565 70.340 205.655 ;
        RECT 71.460 205.225 71.720 205.545 ;
        RECT 72.380 205.225 72.640 205.545 ;
        RECT 71.000 203.525 71.260 203.845 ;
        RECT 70.540 202.505 70.800 202.825 ;
        RECT 69.680 200.895 70.280 201.035 ;
        RECT 67.320 200.125 67.580 200.445 ;
        RECT 68.240 200.125 68.500 200.445 ;
        RECT 69.620 200.125 69.880 200.445 ;
        RECT 67.380 199.280 67.520 200.125 ;
        RECT 67.310 198.910 67.590 199.280 ;
        RECT 68.300 198.345 69.360 198.485 ;
        RECT 68.300 198.065 68.440 198.345 ;
        RECT 66.860 197.745 67.120 198.065 ;
        RECT 68.240 197.745 68.500 198.065 ;
        RECT 66.400 197.065 66.660 197.385 ;
        RECT 68.700 197.065 68.960 197.385 ;
        RECT 68.240 196.385 68.500 196.705 ;
        RECT 68.300 195.345 68.440 196.385 ;
        RECT 68.760 195.345 68.900 197.065 ;
        RECT 68.240 195.025 68.500 195.345 ;
        RECT 68.700 195.025 68.960 195.345 ;
        RECT 69.220 195.005 69.360 198.345 ;
        RECT 69.680 197.385 69.820 200.125 ;
        RECT 69.620 197.065 69.880 197.385 ;
        RECT 70.140 195.200 70.280 200.895 ;
        RECT 70.600 200.445 70.740 202.505 ;
        RECT 71.060 201.885 71.200 203.525 ;
        RECT 71.520 203.165 71.660 205.225 ;
        RECT 71.920 204.545 72.180 204.865 ;
        RECT 71.980 203.165 72.120 204.545 ;
        RECT 72.440 204.040 72.580 205.225 ;
        RECT 72.370 203.670 72.650 204.040 ;
        RECT 71.460 202.845 71.720 203.165 ;
        RECT 71.920 202.845 72.180 203.165 ;
        RECT 71.060 201.745 71.660 201.885 ;
        RECT 71.000 200.805 71.260 201.125 ;
        RECT 71.060 200.445 71.200 200.805 ;
        RECT 70.540 200.125 70.800 200.445 ;
        RECT 71.000 200.125 71.260 200.445 ;
        RECT 66.860 194.685 67.120 195.005 ;
        RECT 67.780 194.685 68.040 195.005 ;
        RECT 69.160 194.685 69.420 195.005 ;
        RECT 70.070 194.830 70.350 195.200 ;
        RECT 65.480 194.405 65.740 194.665 ;
        RECT 66.920 194.405 67.060 194.685 ;
        RECT 67.840 194.520 67.980 194.685 ;
        RECT 65.480 194.345 67.060 194.405 ;
        RECT 63.180 194.005 63.440 194.325 ;
        RECT 65.540 194.265 67.060 194.345 ;
        RECT 63.240 191.945 63.380 194.005 ;
        RECT 62.720 191.625 62.980 191.945 ;
        RECT 63.180 191.625 63.440 191.945 ;
        RECT 62.260 190.945 62.520 191.265 ;
        RECT 64.560 190.945 64.820 191.265 ;
        RECT 62.320 190.245 62.460 190.945 ;
        RECT 62.260 189.925 62.520 190.245 ;
        RECT 64.620 189.610 64.760 190.945 ;
        RECT 66.920 190.245 67.060 194.265 ;
        RECT 67.770 194.150 68.050 194.520 ;
        RECT 70.600 193.985 70.740 200.125 ;
        RECT 70.540 193.665 70.800 193.985 ;
        RECT 70.600 191.945 70.740 193.665 ;
        RECT 71.060 192.965 71.200 200.125 ;
        RECT 71.520 198.405 71.660 201.745 ;
        RECT 72.380 200.125 72.640 200.445 ;
        RECT 71.460 198.085 71.720 198.405 ;
        RECT 71.520 197.725 71.660 198.085 ;
        RECT 72.440 198.065 72.580 200.125 ;
        RECT 72.380 197.745 72.640 198.065 ;
        RECT 71.460 197.405 71.720 197.725 ;
        RECT 72.440 197.385 72.580 197.745 ;
        RECT 71.910 196.870 72.190 197.240 ;
        RECT 72.380 197.065 72.640 197.385 ;
        RECT 71.980 196.705 72.120 196.870 ;
        RECT 72.900 196.705 73.040 213.815 ;
        RECT 74.680 213.725 74.940 214.045 ;
        RECT 73.760 211.005 74.020 211.325 ;
        RECT 74.220 211.005 74.480 211.325 ;
        RECT 73.820 208.945 73.960 211.005 ;
        RECT 74.280 208.945 74.420 211.005 ;
        RECT 74.740 210.160 74.880 213.725 ;
        RECT 75.140 213.385 75.400 213.705 ;
        RECT 75.200 213.025 75.340 213.385 ;
        RECT 75.140 212.705 75.400 213.025 ;
        RECT 75.200 211.665 75.340 212.705 ;
        RECT 75.140 211.345 75.400 211.665 ;
        RECT 76.520 211.235 76.780 211.325 ;
        RECT 76.120 211.095 76.780 211.235 ;
        RECT 76.120 210.895 76.260 211.095 ;
        RECT 76.520 211.005 76.780 211.095 ;
        RECT 75.200 210.755 76.260 210.895 ;
        RECT 74.670 209.790 74.950 210.160 ;
        RECT 73.760 208.625 74.020 208.945 ;
        RECT 74.220 208.625 74.480 208.945 ;
        RECT 73.300 207.265 73.560 207.585 ;
        RECT 73.820 207.495 73.960 208.625 ;
        RECT 74.220 207.495 74.480 207.585 ;
        RECT 73.820 207.355 74.480 207.495 ;
        RECT 74.220 207.265 74.480 207.355 ;
        RECT 73.360 197.725 73.500 207.265 ;
        RECT 74.280 206.225 74.420 207.265 ;
        RECT 74.220 205.905 74.480 206.225 ;
        RECT 73.750 203.670 74.030 204.040 ;
        RECT 73.820 202.825 73.960 203.670 ;
        RECT 74.280 202.825 74.420 205.905 ;
        RECT 73.760 202.505 74.020 202.825 ;
        RECT 74.220 202.505 74.480 202.825 ;
        RECT 73.760 200.465 74.020 200.785 ;
        RECT 73.300 197.405 73.560 197.725 ;
        RECT 73.820 197.045 73.960 200.465 ;
        RECT 74.740 200.105 74.880 209.790 ;
        RECT 75.200 208.265 75.340 210.755 ;
        RECT 76.060 209.985 76.320 210.305 ;
        RECT 76.120 209.480 76.260 209.985 ;
        RECT 75.600 208.965 75.860 209.285 ;
        RECT 76.050 209.110 76.330 209.480 ;
        RECT 77.500 209.285 77.640 216.785 ;
        RECT 78.820 216.105 79.080 216.425 ;
        RECT 79.280 216.105 79.540 216.425 ;
        RECT 77.890 211.830 78.170 212.200 ;
        RECT 78.880 212.005 79.020 216.105 ;
        RECT 79.340 214.920 79.480 216.105 ;
        RECT 79.740 215.765 80.000 216.085 ;
        RECT 79.270 214.550 79.550 214.920 ;
        RECT 79.280 214.405 79.540 214.550 ;
        RECT 79.800 213.365 79.940 215.765 ;
        RECT 81.120 214.405 81.380 214.725 ;
        RECT 79.740 213.045 80.000 213.365 ;
        RECT 81.180 212.005 81.320 214.405 ;
        RECT 77.440 208.965 77.700 209.285 ;
        RECT 75.660 208.265 75.800 208.965 ;
        RECT 76.060 208.625 76.320 208.945 ;
        RECT 75.140 207.945 75.400 208.265 ;
        RECT 75.600 207.945 75.860 208.265 ;
        RECT 74.680 199.785 74.940 200.105 ;
        RECT 74.220 197.405 74.480 197.725 ;
        RECT 74.680 197.405 74.940 197.725 ;
        RECT 73.760 196.725 74.020 197.045 ;
        RECT 71.460 196.385 71.720 196.705 ;
        RECT 71.920 196.385 72.180 196.705 ;
        RECT 72.840 196.385 73.100 196.705 ;
        RECT 73.300 196.560 73.560 196.705 ;
        RECT 71.000 192.645 71.260 192.965 ;
        RECT 69.160 191.625 69.420 191.945 ;
        RECT 70.540 191.625 70.800 191.945 ;
        RECT 66.860 189.925 67.120 190.245 ;
        RECT 69.220 189.610 69.360 191.625 ;
        RECT 71.520 189.905 71.660 196.385 ;
        RECT 71.980 195.880 72.120 196.385 ;
        RECT 73.290 196.190 73.570 196.560 ;
        RECT 71.910 195.510 72.190 195.880 ;
        RECT 74.280 194.665 74.420 197.405 ;
        RECT 74.740 197.240 74.880 197.405 ;
        RECT 74.670 196.870 74.950 197.240 ;
        RECT 74.680 196.385 74.940 196.705 ;
        RECT 74.220 194.345 74.480 194.665 ;
        RECT 72.380 193.665 72.640 193.985 ;
        RECT 74.740 193.840 74.880 196.385 ;
        RECT 71.920 191.855 72.180 191.945 ;
        RECT 72.440 191.855 72.580 193.665 ;
        RECT 74.670 193.470 74.950 193.840 ;
        RECT 75.200 192.965 75.340 207.945 ;
        RECT 76.120 204.865 76.260 208.625 ;
        RECT 76.980 208.285 77.240 208.605 ;
        RECT 76.510 206.390 76.790 206.760 ;
        RECT 76.520 206.245 76.780 206.390 ;
        RECT 76.060 204.775 76.320 204.865 ;
        RECT 75.660 204.635 76.320 204.775 ;
        RECT 75.660 202.825 75.800 204.635 ;
        RECT 76.060 204.545 76.320 204.635 ;
        RECT 77.040 203.845 77.180 208.285 ;
        RECT 76.980 203.525 77.240 203.845 ;
        RECT 75.600 202.505 75.860 202.825 ;
        RECT 76.060 202.505 76.320 202.825 ;
        RECT 76.520 202.505 76.780 202.825 ;
        RECT 76.120 201.125 76.260 202.505 ;
        RECT 76.060 201.035 76.320 201.125 ;
        RECT 75.660 200.895 76.320 201.035 ;
        RECT 75.660 199.425 75.800 200.895 ;
        RECT 76.060 200.805 76.320 200.895 ;
        RECT 76.580 200.785 76.720 202.505 ;
        RECT 76.970 200.950 77.250 201.320 ;
        RECT 76.520 200.465 76.780 200.785 ;
        RECT 77.040 200.445 77.180 200.950 ;
        RECT 76.980 200.125 77.240 200.445 ;
        RECT 77.960 200.105 78.100 211.830 ;
        RECT 78.820 211.685 79.080 212.005 ;
        RECT 81.120 211.685 81.380 212.005 ;
        RECT 82.500 211.685 82.760 212.005 ;
        RECT 79.730 211.150 80.010 211.520 ;
        RECT 82.030 211.150 82.310 211.520 ;
        RECT 78.360 210.665 78.620 210.985 ;
        RECT 78.820 210.840 79.080 210.985 ;
        RECT 78.420 209.285 78.560 210.665 ;
        RECT 78.810 210.470 79.090 210.840 ;
        RECT 78.360 208.965 78.620 209.285 ;
        RECT 78.820 207.945 79.080 208.265 ;
        RECT 78.360 207.605 78.620 207.925 ;
        RECT 77.900 199.785 78.160 200.105 ;
        RECT 75.600 199.105 75.860 199.425 ;
        RECT 77.900 197.295 78.160 197.385 ;
        RECT 78.420 197.295 78.560 207.605 ;
        RECT 78.880 206.565 79.020 207.945 ;
        RECT 79.800 207.925 79.940 211.150 ;
        RECT 82.040 211.005 82.300 211.150 ;
        RECT 80.200 210.325 80.460 210.645 ;
        RECT 81.120 210.325 81.380 210.645 ;
        RECT 79.740 207.605 80.000 207.925 ;
        RECT 79.280 207.265 79.540 207.585 ;
        RECT 78.820 206.245 79.080 206.565 ;
        RECT 78.880 205.545 79.020 206.245 ;
        RECT 79.340 206.225 79.480 207.265 ;
        RECT 79.280 205.905 79.540 206.225 ;
        RECT 78.820 205.225 79.080 205.545 ;
        RECT 78.880 200.445 79.020 205.225 ;
        RECT 78.820 200.125 79.080 200.445 ;
        RECT 79.340 200.015 79.480 205.905 ;
        RECT 79.740 202.505 80.000 202.825 ;
        RECT 79.800 200.785 79.940 202.505 ;
        RECT 79.740 200.465 80.000 200.785 ;
        RECT 79.740 200.015 80.000 200.105 ;
        RECT 79.340 199.875 80.000 200.015 ;
        RECT 80.260 200.015 80.400 210.325 ;
        RECT 81.180 208.265 81.320 210.325 ;
        RECT 82.040 209.985 82.300 210.305 ;
        RECT 80.660 207.945 80.920 208.265 ;
        RECT 81.120 207.945 81.380 208.265 ;
        RECT 80.720 205.545 80.860 207.945 ;
        RECT 81.580 207.605 81.840 207.925 ;
        RECT 81.640 205.885 81.780 207.605 ;
        RECT 82.100 205.885 82.240 209.985 ;
        RECT 81.580 205.565 81.840 205.885 ;
        RECT 82.040 205.565 82.300 205.885 ;
        RECT 80.660 205.225 80.920 205.545 ;
        RECT 81.640 203.845 81.780 205.565 ;
        RECT 81.580 203.525 81.840 203.845 ;
        RECT 82.560 202.565 82.700 211.685 ;
        RECT 82.960 209.985 83.220 210.305 ;
        RECT 83.020 208.605 83.160 209.985 ;
        RECT 82.960 208.285 83.220 208.605 ;
        RECT 83.020 207.440 83.160 208.285 ;
        RECT 83.880 207.945 84.140 208.265 ;
        RECT 82.950 207.070 83.230 207.440 ;
        RECT 83.940 206.565 84.080 207.945 ;
        RECT 83.880 206.245 84.140 206.565 ;
        RECT 84.400 206.225 84.540 218.485 ;
        RECT 86.630 218.265 86.910 219.450 ;
        RECT 98.590 220.190 98.870 221.250 ;
        RECT 110.550 220.945 110.850 221.000 ;
        RECT 110.540 220.600 110.850 220.945 ;
        RECT 98.590 219.790 98.890 220.190 ;
        RECT 86.700 217.885 86.840 218.265 ;
        RECT 98.140 218.145 98.400 218.465 ;
        RECT 98.590 218.265 98.870 219.790 ;
        RECT 99.520 219.505 99.780 219.825 ;
        RECT 86.700 217.745 87.300 217.885 ;
        RECT 84.800 217.125 85.060 217.445 ;
        RECT 84.860 216.425 85.000 217.125 ;
        RECT 84.800 216.105 85.060 216.425 ;
        RECT 84.860 215.745 85.000 216.105 ;
        RECT 87.160 215.745 87.300 217.745 ;
        RECT 91.230 216.590 91.510 216.960 ;
        RECT 84.800 215.425 85.060 215.745 ;
        RECT 86.640 215.425 86.900 215.745 ;
        RECT 87.100 215.425 87.360 215.745 ;
        RECT 85.710 214.550 85.990 214.920 ;
        RECT 85.260 213.045 85.520 213.365 ;
        RECT 85.320 212.005 85.460 213.045 ;
        RECT 85.260 211.685 85.520 212.005 ;
        RECT 85.780 211.405 85.920 214.550 ;
        RECT 86.180 213.725 86.440 214.045 ;
        RECT 86.240 213.560 86.380 213.725 ;
        RECT 86.170 213.190 86.450 213.560 ;
        RECT 86.700 212.005 86.840 215.425 ;
        RECT 90.310 213.870 90.590 214.240 ;
        RECT 87.090 213.190 87.370 213.560 ;
        RECT 88.480 213.385 88.740 213.705 ;
        RECT 86.640 211.685 86.900 212.005 ;
        RECT 84.800 211.005 85.060 211.325 ;
        RECT 85.780 211.265 86.840 211.405 ;
        RECT 87.160 211.325 87.300 213.190 ;
        RECT 84.860 210.305 85.000 211.005 ;
        RECT 84.800 209.985 85.060 210.305 ;
        RECT 85.780 208.605 85.920 211.265 ;
        RECT 86.180 210.665 86.440 210.985 ;
        RECT 86.700 210.725 86.840 211.265 ;
        RECT 87.100 211.005 87.360 211.325 ;
        RECT 87.560 211.005 87.820 211.325 ;
        RECT 87.620 210.725 87.760 211.005 ;
        RECT 88.540 210.985 88.680 213.385 ;
        RECT 89.860 213.045 90.120 213.365 ;
        RECT 89.920 212.005 90.060 213.045 ;
        RECT 89.860 211.685 90.120 212.005 ;
        RECT 86.240 209.285 86.380 210.665 ;
        RECT 86.700 210.585 87.760 210.725 ;
        RECT 88.480 210.665 88.740 210.985 ;
        RECT 88.940 210.325 89.200 210.645 ;
        RECT 86.640 209.985 86.900 210.305 ;
        RECT 86.180 208.965 86.440 209.285 ;
        RECT 85.720 208.515 85.980 208.605 ;
        RECT 85.320 208.375 85.980 208.515 ;
        RECT 84.340 205.905 84.600 206.225 ;
        RECT 83.880 204.545 84.140 204.865 ;
        RECT 83.940 203.165 84.080 204.545 ;
        RECT 83.880 202.845 84.140 203.165 ;
        RECT 84.800 202.845 85.060 203.165 ;
        RECT 82.100 202.425 82.700 202.565 ;
        RECT 83.420 202.505 83.680 202.825 ;
        RECT 81.120 200.125 81.380 200.445 ;
        RECT 80.660 200.015 80.920 200.105 ;
        RECT 80.260 199.875 80.920 200.015 ;
        RECT 78.820 199.105 79.080 199.425 ;
        RECT 78.880 197.385 79.020 199.105 ;
        RECT 77.900 197.155 78.560 197.295 ;
        RECT 77.900 197.065 78.160 197.155 ;
        RECT 78.820 197.065 79.080 197.385 ;
        RECT 76.520 196.385 76.780 196.705 ;
        RECT 76.580 195.255 76.720 196.385 ;
        RECT 76.980 195.255 77.240 195.345 ;
        RECT 76.580 195.115 77.240 195.255 ;
        RECT 76.980 195.025 77.240 195.115 ;
        RECT 75.140 192.645 75.400 192.965 ;
        RECT 77.040 192.625 77.180 195.025 ;
        RECT 78.820 194.345 79.080 194.665 ;
        RECT 76.980 192.305 77.240 192.625 ;
        RECT 78.880 191.945 79.020 194.345 ;
        RECT 79.340 192.285 79.480 199.875 ;
        RECT 79.740 199.785 80.000 199.875 ;
        RECT 80.660 199.785 80.920 199.875 ;
        RECT 80.200 199.105 80.460 199.425 ;
        RECT 79.740 196.725 80.000 197.045 ;
        RECT 79.800 192.965 79.940 196.725 ;
        RECT 80.260 195.005 80.400 199.105 ;
        RECT 80.660 197.065 80.920 197.385 ;
        RECT 80.720 195.685 80.860 197.065 ;
        RECT 80.660 195.365 80.920 195.685 ;
        RECT 81.180 195.345 81.320 200.125 ;
        RECT 81.570 196.870 81.850 197.240 ;
        RECT 81.640 196.705 81.780 196.870 ;
        RECT 81.580 196.385 81.840 196.705 ;
        RECT 82.100 195.345 82.240 202.425 ;
        RECT 82.500 201.825 82.760 202.145 ;
        RECT 81.120 195.025 81.380 195.345 ;
        RECT 82.040 195.025 82.300 195.345 ;
        RECT 82.560 195.200 82.700 201.825 ;
        RECT 83.480 200.785 83.620 202.505 ;
        RECT 84.860 202.145 85.000 202.845 ;
        RECT 85.320 202.825 85.460 208.375 ;
        RECT 85.720 208.285 85.980 208.375 ;
        RECT 86.180 207.265 86.440 207.585 ;
        RECT 86.240 205.885 86.380 207.265 ;
        RECT 86.700 205.885 86.840 209.985 ;
        RECT 87.100 208.285 87.360 208.605 ;
        RECT 87.160 207.440 87.300 208.285 ;
        RECT 87.560 207.945 87.820 208.265 ;
        RECT 88.020 207.945 88.280 208.265 ;
        RECT 88.480 208.175 88.740 208.265 ;
        RECT 89.000 208.175 89.140 210.325 ;
        RECT 88.480 208.035 90.060 208.175 ;
        RECT 88.480 207.945 88.740 208.035 ;
        RECT 87.090 207.070 87.370 207.440 ;
        RECT 87.620 206.225 87.760 207.945 ;
        RECT 87.560 205.905 87.820 206.225 ;
        RECT 86.180 205.565 86.440 205.885 ;
        RECT 86.640 205.565 86.900 205.885 ;
        RECT 88.080 205.545 88.220 207.945 ;
        RECT 89.390 205.710 89.670 206.080 ;
        RECT 85.720 204.885 85.980 205.205 ;
        RECT 86.630 205.030 86.910 205.400 ;
        RECT 88.020 205.225 88.280 205.545 ;
        RECT 86.640 204.885 86.900 205.030 ;
        RECT 85.260 202.505 85.520 202.825 ;
        RECT 84.800 201.825 85.060 202.145 ;
        RECT 83.420 200.465 83.680 200.785 ;
        RECT 84.340 200.465 84.600 200.785 ;
        RECT 82.960 199.445 83.220 199.765 ;
        RECT 83.020 199.280 83.160 199.445 ;
        RECT 82.950 198.910 83.230 199.280 ;
        RECT 83.020 195.880 83.160 198.910 ;
        RECT 83.480 198.405 83.620 200.465 ;
        RECT 83.880 199.785 84.140 200.105 ;
        RECT 83.420 198.085 83.680 198.405 ;
        RECT 83.940 196.615 84.080 199.785 ;
        RECT 84.400 197.385 84.540 200.465 ;
        RECT 84.860 197.385 85.000 201.825 ;
        RECT 85.320 200.445 85.460 202.505 ;
        RECT 85.260 200.125 85.520 200.445 ;
        RECT 85.780 199.845 85.920 204.885 ;
        RECT 87.090 204.350 87.370 204.720 ;
        RECT 88.940 204.545 89.200 204.865 ;
        RECT 87.160 203.165 87.300 204.350 ;
        RECT 88.020 203.525 88.280 203.845 ;
        RECT 87.560 203.360 87.820 203.505 ;
        RECT 87.100 202.845 87.360 203.165 ;
        RECT 87.550 202.990 87.830 203.360 ;
        RECT 88.080 202.565 88.220 203.525 ;
        RECT 89.000 203.505 89.140 204.545 ;
        RECT 88.940 203.185 89.200 203.505 ;
        RECT 89.460 202.825 89.600 205.710 ;
        RECT 88.940 202.565 89.200 202.825 ;
        RECT 88.080 202.505 89.200 202.565 ;
        RECT 89.400 202.505 89.660 202.825 ;
        RECT 88.080 202.425 89.140 202.505 ;
        RECT 88.080 200.445 88.220 202.425 ;
        RECT 88.940 201.825 89.200 202.145 ;
        RECT 89.400 202.000 89.660 202.145 ;
        RECT 89.000 200.445 89.140 201.825 ;
        RECT 89.390 201.630 89.670 202.000 ;
        RECT 89.920 201.205 90.060 208.035 ;
        RECT 90.380 205.205 90.520 213.870 ;
        RECT 91.300 211.665 91.440 216.590 ;
        RECT 97.220 216.445 97.480 216.765 ;
        RECT 94.460 215.425 94.720 215.745 ;
        RECT 91.690 214.550 91.970 214.920 ;
        RECT 91.240 211.345 91.500 211.665 ;
        RECT 90.780 211.005 91.040 211.325 ;
        RECT 90.840 210.305 90.980 211.005 ;
        RECT 90.780 209.985 91.040 210.305 ;
        RECT 90.840 208.945 90.980 209.985 ;
        RECT 90.780 208.625 91.040 208.945 ;
        RECT 90.840 205.545 90.980 208.625 ;
        RECT 91.240 207.945 91.500 208.265 ;
        RECT 91.300 206.225 91.440 207.945 ;
        RECT 91.240 205.905 91.500 206.225 ;
        RECT 90.780 205.225 91.040 205.545 ;
        RECT 90.320 204.885 90.580 205.205 ;
        RECT 90.840 204.605 90.980 205.225 ;
        RECT 89.460 201.065 90.060 201.205 ;
        RECT 90.380 204.465 90.980 204.605 ;
        RECT 88.020 200.125 88.280 200.445 ;
        RECT 88.940 200.125 89.200 200.445 ;
        RECT 85.320 199.705 85.920 199.845 ;
        RECT 84.340 197.065 84.600 197.385 ;
        RECT 84.800 197.065 85.060 197.385 ;
        RECT 84.860 196.615 85.000 197.065 ;
        RECT 83.940 196.475 85.000 196.615 ;
        RECT 82.950 195.510 83.230 195.880 ;
        RECT 80.200 194.685 80.460 195.005 ;
        RECT 82.490 194.830 82.770 195.200 ;
        RECT 79.740 192.645 80.000 192.965 ;
        RECT 79.280 191.965 79.540 192.285 ;
        RECT 80.260 191.945 80.400 194.685 ;
        RECT 82.960 193.665 83.220 193.985 ;
        RECT 83.020 191.945 83.160 193.665 ;
        RECT 83.940 192.625 84.080 196.475 ;
        RECT 85.320 195.685 85.460 199.705 ;
        RECT 86.180 199.105 86.440 199.425 ;
        RECT 87.100 199.280 87.360 199.425 ;
        RECT 86.240 197.725 86.380 199.105 ;
        RECT 87.090 198.910 87.370 199.280 ;
        RECT 86.180 197.405 86.440 197.725 ;
        RECT 85.260 195.365 85.520 195.685 ;
        RECT 84.800 194.345 85.060 194.665 ;
        RECT 84.860 192.965 85.000 194.345 ;
        RECT 86.240 192.965 86.380 197.405 ;
        RECT 88.020 196.725 88.280 197.045 ;
        RECT 88.080 195.685 88.220 196.725 ;
        RECT 88.020 195.365 88.280 195.685 ;
        RECT 84.800 192.645 85.060 192.965 ;
        RECT 86.180 192.645 86.440 192.965 ;
        RECT 83.880 192.305 84.140 192.625 ;
        RECT 88.080 191.945 88.220 195.365 ;
        RECT 89.460 191.945 89.600 201.065 ;
        RECT 90.380 200.785 90.520 204.465 ;
        RECT 91.760 202.825 91.900 214.550 ;
        RECT 94.520 211.325 94.660 215.425 ;
        RECT 97.280 214.725 97.420 216.445 ;
        RECT 98.200 216.085 98.340 218.145 ;
        RECT 98.660 216.765 98.800 218.265 ;
        RECT 98.600 216.445 98.860 216.765 ;
        RECT 99.060 216.105 99.320 216.425 ;
        RECT 97.680 215.765 97.940 216.085 ;
        RECT 98.140 215.765 98.400 216.085 ;
        RECT 97.220 214.405 97.480 214.725 ;
        RECT 97.740 214.240 97.880 215.765 ;
        RECT 97.670 213.870 97.950 214.240 ;
        RECT 97.210 211.830 97.490 212.200 ;
        RECT 97.280 211.665 97.420 211.830 ;
        RECT 96.760 211.345 97.020 211.665 ;
        RECT 97.220 211.345 97.480 211.665 ;
        RECT 93.080 211.005 93.340 211.325 ;
        RECT 94.460 211.005 94.720 211.325 ;
        RECT 93.140 209.285 93.280 211.005 ;
        RECT 94.000 209.985 94.260 210.305 ;
        RECT 93.080 208.965 93.340 209.285 ;
        RECT 94.060 207.925 94.200 209.985 ;
        RECT 95.840 208.625 96.100 208.945 ;
        RECT 94.920 208.175 95.180 208.265 ;
        RECT 95.900 208.175 96.040 208.625 ;
        RECT 96.290 208.430 96.570 208.800 ;
        RECT 94.920 208.035 96.040 208.175 ;
        RECT 94.920 207.945 95.180 208.035 ;
        RECT 92.620 207.605 92.880 207.925 ;
        RECT 94.000 207.605 94.260 207.925 ;
        RECT 94.460 207.605 94.720 207.925 ;
        RECT 92.680 205.885 92.820 207.605 ;
        RECT 93.540 207.440 93.800 207.585 ;
        RECT 93.530 207.325 93.810 207.440 ;
        RECT 93.140 207.185 93.810 207.325 ;
        RECT 92.620 205.565 92.880 205.885 ;
        RECT 92.680 204.865 92.820 205.565 ;
        RECT 92.620 204.545 92.880 204.865 ;
        RECT 91.700 202.505 91.960 202.825 ;
        RECT 92.150 202.310 92.430 202.680 ;
        RECT 92.220 202.145 92.360 202.310 ;
        RECT 90.780 201.825 91.040 202.145 ;
        RECT 92.160 201.825 92.420 202.145 ;
        RECT 90.320 200.465 90.580 200.785 ;
        RECT 90.840 200.640 90.980 201.825 ;
        RECT 93.140 200.640 93.280 207.185 ;
        RECT 93.530 207.070 93.810 207.185 ;
        RECT 94.520 205.885 94.660 207.605 ;
        RECT 94.460 205.565 94.720 205.885 ;
        RECT 93.530 202.990 93.810 203.360 ;
        RECT 93.600 202.825 93.740 202.990 ;
        RECT 94.000 202.845 94.260 203.165 ;
        RECT 93.540 202.505 93.800 202.825 ;
        RECT 94.060 202.680 94.200 202.845 ;
        RECT 93.990 202.310 94.270 202.680 ;
        RECT 93.540 201.825 93.800 202.145 ;
        RECT 90.770 200.270 91.050 200.640 ;
        RECT 93.070 200.525 93.350 200.640 ;
        RECT 92.680 200.445 93.350 200.525 ;
        RECT 92.620 200.385 93.350 200.445 ;
        RECT 92.620 200.125 92.880 200.385 ;
        RECT 93.070 200.270 93.350 200.385 ;
        RECT 93.080 199.785 93.340 200.105 ;
        RECT 91.700 197.065 91.960 197.385 ;
        RECT 89.860 196.725 90.120 197.045 ;
        RECT 71.920 191.715 72.580 191.855 ;
        RECT 71.920 191.625 72.180 191.715 ;
        RECT 78.820 191.625 79.080 191.945 ;
        RECT 80.200 191.625 80.460 191.945 ;
        RECT 82.960 191.625 83.220 191.945 ;
        RECT 87.100 191.855 87.360 191.945 ;
        RECT 87.100 191.715 87.760 191.855 ;
        RECT 87.100 191.625 87.360 191.715 ;
        RECT 78.360 191.285 78.620 191.605 ;
        RECT 79.740 191.285 80.000 191.605 ;
        RECT 73.760 190.945 74.020 191.265 ;
        RECT 73.820 190.060 73.960 190.945 ;
        RECT 78.420 190.060 78.560 191.285 ;
        RECT 79.800 190.245 79.940 191.285 ;
        RECT 82.960 190.945 83.220 191.265 ;
        RECT 73.820 189.920 78.560 190.060 ;
        RECT 79.740 189.925 80.000 190.245 ;
        RECT 64.620 189.470 69.360 189.610 ;
        RECT 71.460 189.585 71.720 189.905 ;
        RECT 61.800 188.905 62.060 189.225 ;
        RECT 60.420 187.885 60.680 188.205 ;
        RECT 64.620 187.715 64.760 189.470 ;
        RECT 69.220 187.715 69.360 189.470 ;
        RECT 73.820 187.715 73.960 189.920 ;
        RECT 78.420 187.715 78.560 189.920 ;
        RECT 83.020 189.910 83.160 190.945 ;
        RECT 87.620 189.910 87.760 191.715 ;
        RECT 88.020 191.625 88.280 191.945 ;
        RECT 89.400 191.625 89.660 191.945 ;
        RECT 88.480 191.285 88.740 191.605 ;
        RECT 88.540 190.245 88.680 191.285 ;
        RECT 89.460 191.265 89.600 191.625 ;
        RECT 89.920 191.605 90.060 196.725 ;
        RECT 91.760 193.985 91.900 197.065 ;
        RECT 93.140 197.045 93.280 199.785 ;
        RECT 93.080 196.725 93.340 197.045 ;
        RECT 92.620 196.385 92.880 196.705 ;
        RECT 91.700 193.665 91.960 193.985 ;
        RECT 92.680 191.945 92.820 196.385 ;
        RECT 93.080 194.345 93.340 194.665 ;
        RECT 93.140 192.965 93.280 194.345 ;
        RECT 93.080 192.645 93.340 192.965 ;
        RECT 92.620 191.625 92.880 191.945 ;
        RECT 89.860 191.285 90.120 191.605 ;
        RECT 89.400 190.945 89.660 191.265 ;
        RECT 92.160 190.945 92.420 191.265 ;
        RECT 88.480 189.925 88.740 190.245 ;
        RECT 83.020 189.770 87.760 189.910 ;
        RECT 83.020 187.715 83.160 189.770 ;
        RECT 87.620 187.715 87.760 189.770 ;
        RECT 89.460 189.225 89.600 190.945 ;
        RECT 89.400 188.905 89.660 189.225 ;
        RECT 92.220 187.715 92.360 190.945 ;
        RECT 93.600 187.825 93.740 201.825 ;
        RECT 94.520 199.425 94.660 205.565 ;
        RECT 94.980 200.445 95.120 207.945 ;
        RECT 96.360 207.925 96.500 208.430 ;
        RECT 96.300 207.605 96.560 207.925 ;
        RECT 96.360 202.825 96.500 207.605 ;
        RECT 96.820 205.885 96.960 211.345 ;
        RECT 97.740 208.265 97.880 213.870 ;
        RECT 98.140 212.705 98.400 213.025 ;
        RECT 98.200 210.645 98.340 212.705 ;
        RECT 98.600 211.685 98.860 212.005 ;
        RECT 98.140 210.325 98.400 210.645 ;
        RECT 98.660 209.365 98.800 211.685 ;
        RECT 98.200 209.225 98.800 209.365 ;
        RECT 97.680 207.945 97.940 208.265 ;
        RECT 97.740 207.440 97.880 207.945 ;
        RECT 97.670 207.070 97.950 207.440 ;
        RECT 96.760 205.565 97.020 205.885 ;
        RECT 96.820 203.505 96.960 205.565 ;
        RECT 97.680 204.885 97.940 205.205 ;
        RECT 96.760 203.185 97.020 203.505 ;
        RECT 96.300 202.505 96.560 202.825 ;
        RECT 95.840 200.465 96.100 200.785 ;
        RECT 94.920 200.125 95.180 200.445 ;
        RECT 94.460 199.105 94.720 199.425 ;
        RECT 94.520 192.625 94.660 199.105 ;
        RECT 95.370 198.230 95.650 198.600 ;
        RECT 95.440 197.725 95.580 198.230 ;
        RECT 95.380 197.405 95.640 197.725 ;
        RECT 94.460 192.305 94.720 192.625 ;
        RECT 95.900 192.285 96.040 200.465 ;
        RECT 96.360 197.385 96.500 202.505 ;
        RECT 96.820 200.445 96.960 203.185 ;
        RECT 97.740 202.825 97.880 204.885 ;
        RECT 97.220 202.505 97.480 202.825 ;
        RECT 97.680 202.505 97.940 202.825 ;
        RECT 97.280 202.145 97.420 202.505 ;
        RECT 97.220 201.825 97.480 202.145 ;
        RECT 97.280 201.320 97.420 201.825 ;
        RECT 97.210 200.950 97.490 201.320 ;
        RECT 97.740 201.125 97.880 202.505 ;
        RECT 98.200 201.320 98.340 209.225 ;
        RECT 98.600 208.685 98.860 208.945 ;
        RECT 99.120 208.685 99.260 216.105 ;
        RECT 99.580 216.085 99.720 219.505 ;
        RECT 110.540 219.340 110.830 220.600 ;
        RECT 103.200 218.145 103.460 218.465 ;
        RECT 110.550 218.265 110.830 219.340 ;
        RECT 122.510 218.265 122.790 221.900 ;
        RECT 133.560 218.825 133.820 219.145 ;
        RECT 102.740 216.105 103.000 216.425 ;
        RECT 99.520 215.765 99.780 216.085 ;
        RECT 100.440 215.425 100.700 215.745 ;
        RECT 99.980 214.065 100.240 214.385 ;
        RECT 100.040 211.665 100.180 214.065 ;
        RECT 99.980 211.345 100.240 211.665 ;
        RECT 98.600 208.625 99.260 208.685 ;
        RECT 98.660 208.545 99.260 208.625 ;
        RECT 99.120 208.265 99.260 208.545 ;
        RECT 99.980 208.285 100.240 208.605 ;
        RECT 99.060 207.945 99.320 208.265 ;
        RECT 99.520 207.945 99.780 208.265 ;
        RECT 99.580 207.585 99.720 207.945 ;
        RECT 99.520 207.265 99.780 207.585 ;
        RECT 99.060 206.475 99.320 206.565 ;
        RECT 100.040 206.475 100.180 208.285 ;
        RECT 99.060 206.335 100.180 206.475 ;
        RECT 99.060 206.245 99.320 206.335 ;
        RECT 98.600 205.225 98.860 205.545 ;
        RECT 98.660 202.825 98.800 205.225 ;
        RECT 98.600 202.505 98.860 202.825 ;
        RECT 97.680 200.805 97.940 201.125 ;
        RECT 98.130 200.950 98.410 201.320 ;
        RECT 98.140 200.805 98.400 200.950 ;
        RECT 99.120 200.445 99.260 206.245 ;
        RECT 99.520 204.885 99.780 205.205 ;
        RECT 99.580 203.505 99.720 204.885 ;
        RECT 99.520 203.185 99.780 203.505 ;
        RECT 100.500 202.825 100.640 215.425 ;
        RECT 102.800 214.385 102.940 216.105 ;
        RECT 102.740 214.065 103.000 214.385 ;
        RECT 101.360 213.725 101.620 214.045 ;
        RECT 100.900 213.385 101.160 213.705 ;
        RECT 100.960 208.945 101.100 213.385 ;
        RECT 100.900 208.625 101.160 208.945 ;
        RECT 100.890 207.750 101.170 208.120 ;
        RECT 100.960 205.885 101.100 207.750 ;
        RECT 100.900 205.565 101.160 205.885 ;
        RECT 101.420 203.165 101.560 213.725 ;
        RECT 101.820 213.560 102.080 213.705 ;
        RECT 101.810 213.190 102.090 213.560 ;
        RECT 102.270 212.510 102.550 212.880 ;
        RECT 102.340 210.215 102.480 212.510 ;
        RECT 101.880 210.075 102.480 210.215 ;
        RECT 101.360 202.845 101.620 203.165 ;
        RECT 99.520 202.505 99.780 202.825 ;
        RECT 100.440 202.505 100.700 202.825 ;
        RECT 99.580 201.125 99.720 202.505 ;
        RECT 100.500 202.145 100.640 202.505 ;
        RECT 101.350 202.310 101.630 202.680 ;
        RECT 101.420 202.145 101.560 202.310 ;
        RECT 100.440 201.825 100.700 202.145 ;
        RECT 101.360 201.825 101.620 202.145 ;
        RECT 99.520 200.805 99.780 201.125 ;
        RECT 96.760 200.125 97.020 200.445 ;
        RECT 99.060 200.125 99.320 200.445 ;
        RECT 99.580 199.845 99.720 200.805 ;
        RECT 100.440 200.465 100.700 200.785 ;
        RECT 100.500 200.105 100.640 200.465 ;
        RECT 101.420 200.105 101.560 201.825 ;
        RECT 101.880 200.445 102.020 210.075 ;
        RECT 102.280 207.945 102.540 208.265 ;
        RECT 102.340 202.825 102.480 207.945 ;
        RECT 102.730 206.390 103.010 206.760 ;
        RECT 102.740 206.245 103.000 206.390 ;
        RECT 103.260 203.925 103.400 218.145 ;
        RECT 110.620 218.065 110.760 218.265 ;
        RECT 122.575 218.045 122.715 218.265 ;
        RECT 122.575 217.905 125.480 218.045 ;
        RECT 105.500 217.125 105.760 217.445 ;
        RECT 103.660 216.785 103.920 217.105 ;
        RECT 103.720 207.925 103.860 216.785 ;
        RECT 104.120 213.045 104.380 213.365 ;
        RECT 104.180 212.005 104.320 213.045 ;
        RECT 105.040 212.705 105.300 213.025 ;
        RECT 105.100 212.005 105.240 212.705 ;
        RECT 104.120 211.685 104.380 212.005 ;
        RECT 105.040 211.685 105.300 212.005 ;
        RECT 104.180 208.605 104.320 211.685 ;
        RECT 105.560 211.325 105.700 217.125 ;
        RECT 125.340 216.845 125.480 217.905 ;
        RECT 125.740 216.845 126.000 217.105 ;
        RECT 125.340 216.785 126.000 216.845 ;
        RECT 124.820 216.445 125.080 216.765 ;
        RECT 125.340 216.705 125.940 216.785 ;
        RECT 127.580 216.445 127.840 216.765 ;
        RECT 128.500 216.445 128.760 216.765 ;
        RECT 107.340 216.335 107.600 216.425 ;
        RECT 107.340 216.195 108.000 216.335 ;
        RECT 107.340 216.105 107.600 216.195 ;
        RECT 106.420 213.385 106.680 213.705 ;
        RECT 106.880 213.385 107.140 213.705 ;
        RECT 105.960 212.705 106.220 213.025 ;
        RECT 105.500 211.005 105.760 211.325 ;
        RECT 104.120 208.515 104.380 208.605 ;
        RECT 104.120 208.375 104.780 208.515 ;
        RECT 105.030 208.430 105.310 208.800 ;
        RECT 104.120 208.285 104.380 208.375 ;
        RECT 103.660 207.605 103.920 207.925 ;
        RECT 104.120 207.265 104.380 207.585 ;
        RECT 103.650 206.390 103.930 206.760 ;
        RECT 103.720 204.865 103.860 206.390 ;
        RECT 104.180 205.885 104.320 207.265 ;
        RECT 104.640 205.885 104.780 208.375 ;
        RECT 105.100 208.265 105.240 208.430 ;
        RECT 105.040 207.945 105.300 208.265 ;
        RECT 105.100 207.585 105.240 207.945 ;
        RECT 105.040 207.265 105.300 207.585 ;
        RECT 105.560 207.440 105.700 211.005 ;
        RECT 105.490 207.070 105.770 207.440 ;
        RECT 106.020 206.225 106.160 212.705 ;
        RECT 106.480 208.800 106.620 213.385 ;
        RECT 106.940 209.285 107.080 213.385 ;
        RECT 107.860 210.645 108.000 216.195 ;
        RECT 108.720 216.105 108.980 216.425 ;
        RECT 112.400 216.105 112.660 216.425 ;
        RECT 108.780 214.725 108.920 216.105 ;
        RECT 108.720 214.405 108.980 214.725 ;
        RECT 108.720 213.385 108.980 213.705 ;
        RECT 108.260 213.045 108.520 213.365 ;
        RECT 108.320 212.200 108.460 213.045 ;
        RECT 108.250 211.830 108.530 212.200 ;
        RECT 108.260 211.005 108.520 211.325 ;
        RECT 107.800 210.325 108.060 210.645 ;
        RECT 106.880 208.965 107.140 209.285 ;
        RECT 106.410 208.430 106.690 208.800 ;
        RECT 105.500 205.905 105.760 206.225 ;
        RECT 105.960 205.905 106.220 206.225 ;
        RECT 104.120 205.565 104.380 205.885 ;
        RECT 104.580 205.565 104.840 205.885 ;
        RECT 105.040 204.885 105.300 205.205 ;
        RECT 103.660 204.545 103.920 204.865 ;
        RECT 102.800 203.785 103.400 203.925 ;
        RECT 102.280 202.505 102.540 202.825 ;
        RECT 102.340 200.785 102.480 202.505 ;
        RECT 102.800 202.145 102.940 203.785 ;
        RECT 103.190 202.310 103.470 202.680 ;
        RECT 102.740 201.825 103.000 202.145 ;
        RECT 102.730 200.950 103.010 201.320 ;
        RECT 102.280 200.465 102.540 200.785 ;
        RECT 101.820 200.125 102.080 200.445 ;
        RECT 96.760 199.445 97.020 199.765 ;
        RECT 97.740 199.705 99.720 199.845 ;
        RECT 100.440 199.785 100.700 200.105 ;
        RECT 101.360 199.785 101.620 200.105 ;
        RECT 102.800 200.015 102.940 200.950 ;
        RECT 103.260 200.445 103.400 202.310 ;
        RECT 103.720 202.145 103.860 204.545 ;
        RECT 104.120 203.185 104.380 203.505 ;
        RECT 104.180 202.680 104.320 203.185 ;
        RECT 104.110 202.310 104.390 202.680 ;
        RECT 104.580 202.505 104.840 202.825 ;
        RECT 103.660 201.825 103.920 202.145 ;
        RECT 104.120 201.825 104.380 202.145 ;
        RECT 103.660 200.465 103.920 200.785 ;
        RECT 103.200 200.125 103.460 200.445 ;
        RECT 102.340 199.875 102.940 200.015 ;
        RECT 96.300 197.065 96.560 197.385 ;
        RECT 96.820 197.295 96.960 199.445 ;
        RECT 97.740 198.405 97.880 199.705 ;
        RECT 99.060 199.105 99.320 199.425 ;
        RECT 100.900 199.165 101.160 199.425 ;
        RECT 100.900 199.105 101.560 199.165 ;
        RECT 97.680 198.085 97.940 198.405 ;
        RECT 97.220 197.805 97.480 198.065 ;
        RECT 98.600 197.805 98.860 198.065 ;
        RECT 97.220 197.745 98.860 197.805 ;
        RECT 99.120 197.805 99.260 199.105 ;
        RECT 100.960 199.025 101.560 199.105 ;
        RECT 101.420 198.600 101.560 199.025 ;
        RECT 100.430 198.230 100.710 198.600 ;
        RECT 101.350 198.230 101.630 198.600 ;
        RECT 97.280 197.665 98.800 197.745 ;
        RECT 99.120 197.665 99.720 197.805 ;
        RECT 100.500 197.725 100.640 198.230 ;
        RECT 96.820 197.155 97.420 197.295 ;
        RECT 96.760 194.345 97.020 194.665 ;
        RECT 95.840 191.965 96.100 192.285 ;
        RECT 94.000 190.945 94.260 191.265 ;
        RECT 94.060 190.245 94.200 190.945 ;
        RECT 94.000 189.925 94.260 190.245 ;
        RECT 13.950 187.290 14.230 187.715 ;
        RECT 18.550 187.290 18.830 187.715 ;
        RECT 23.150 187.590 23.430 187.715 ;
        RECT 13.940 186.890 14.240 187.290 ;
        RECT 18.540 186.890 18.840 187.290 ;
        RECT 23.140 187.190 23.440 187.590 ;
        RECT 13.950 185.715 14.230 186.890 ;
        RECT 18.550 185.715 18.830 186.890 ;
        RECT 23.150 185.715 23.430 187.190 ;
        RECT 27.750 185.715 28.030 187.715 ;
        RECT 32.350 185.840 32.630 187.715 ;
        RECT 32.340 185.440 32.640 185.840 ;
        RECT 36.950 185.715 37.230 187.715 ;
        RECT 41.550 185.715 41.830 187.715 ;
        RECT 46.150 185.715 46.430 187.715 ;
        RECT 50.750 185.715 51.030 187.715 ;
        RECT 55.350 187.510 55.630 187.715 ;
        RECT 59.950 187.510 60.230 187.715 ;
        RECT 55.350 187.370 60.230 187.510 ;
        RECT 55.350 185.715 55.630 187.370 ;
        RECT 59.950 185.715 60.230 187.370 ;
        RECT 64.550 185.715 64.830 187.715 ;
        RECT 69.150 185.715 69.430 187.715 ;
        RECT 73.750 185.715 74.030 187.715 ;
        RECT 78.350 185.715 78.630 187.715 ;
        RECT 82.950 185.715 83.230 187.715 ;
        RECT 87.550 185.715 87.830 187.715 ;
        RECT 92.150 187.160 92.430 187.715 ;
        RECT 93.540 187.505 93.800 187.825 ;
        RECT 96.820 187.715 96.960 194.345 ;
        RECT 97.280 192.965 97.420 197.155 ;
        RECT 99.580 197.045 99.720 197.665 ;
        RECT 100.440 197.405 100.700 197.725 ;
        RECT 102.340 197.385 102.480 199.875 ;
        RECT 103.720 199.675 103.860 200.465 ;
        RECT 104.180 200.445 104.320 201.825 ;
        RECT 104.640 200.445 104.780 202.505 ;
        RECT 105.100 201.125 105.240 204.885 ;
        RECT 105.560 202.145 105.700 205.905 ;
        RECT 105.500 201.825 105.760 202.145 ;
        RECT 105.040 200.805 105.300 201.125 ;
        RECT 105.560 200.445 105.700 201.825 ;
        RECT 104.120 200.125 104.380 200.445 ;
        RECT 104.580 200.125 104.840 200.445 ;
        RECT 105.500 200.125 105.760 200.445 ;
        RECT 105.040 199.675 105.300 199.765 ;
        RECT 103.720 199.535 105.300 199.675 ;
        RECT 105.040 199.445 105.300 199.535 ;
        RECT 102.740 199.105 103.000 199.425 ;
        RECT 102.800 197.920 102.940 199.105 ;
        RECT 105.560 198.405 105.700 200.125 ;
        RECT 105.500 198.085 105.760 198.405 ;
        RECT 106.480 198.065 106.620 208.430 ;
        RECT 107.860 208.265 108.000 210.325 ;
        RECT 107.800 207.945 108.060 208.265 ;
        RECT 108.320 206.565 108.460 211.005 ;
        RECT 108.260 206.245 108.520 206.565 ;
        RECT 107.340 205.225 107.600 205.545 ;
        RECT 107.400 203.845 107.540 205.225 ;
        RECT 107.800 204.885 108.060 205.205 ;
        RECT 106.880 203.525 107.140 203.845 ;
        RECT 107.340 203.525 107.600 203.845 ;
        RECT 106.940 202.825 107.080 203.525 ;
        RECT 107.860 203.165 108.000 204.885 ;
        RECT 107.800 202.845 108.060 203.165 ;
        RECT 106.880 202.680 107.140 202.825 ;
        RECT 106.870 202.310 107.150 202.680 ;
        RECT 107.800 200.695 108.060 200.785 ;
        RECT 108.320 200.695 108.460 206.245 ;
        RECT 107.800 200.555 108.460 200.695 ;
        RECT 107.800 200.465 108.060 200.555 ;
        RECT 107.340 199.105 107.600 199.425 ;
        RECT 102.730 197.550 103.010 197.920 ;
        RECT 104.120 197.745 104.380 198.065 ;
        RECT 104.580 197.745 104.840 198.065 ;
        RECT 106.420 197.745 106.680 198.065 ;
        RECT 104.180 197.385 104.320 197.745 ;
        RECT 102.280 197.065 102.540 197.385 ;
        RECT 102.740 197.065 103.000 197.385 ;
        RECT 104.120 197.065 104.380 197.385 ;
        RECT 99.060 196.725 99.320 197.045 ;
        RECT 99.520 196.725 99.780 197.045 ;
        RECT 98.600 194.685 98.860 195.005 ;
        RECT 98.660 194.325 98.800 194.685 ;
        RECT 98.600 194.005 98.860 194.325 ;
        RECT 97.220 192.645 97.480 192.965 ;
        RECT 97.680 192.305 97.940 192.625 ;
        RECT 97.740 191.945 97.880 192.305 ;
        RECT 97.680 191.625 97.940 191.945 ;
        RECT 99.120 191.605 99.260 196.725 ;
        RECT 99.580 195.345 99.720 196.725 ;
        RECT 99.980 196.385 100.240 196.705 ;
        RECT 100.440 196.385 100.700 196.705 ;
        RECT 99.520 195.025 99.780 195.345 ;
        RECT 100.040 194.665 100.180 196.385 ;
        RECT 99.980 194.345 100.240 194.665 ;
        RECT 100.500 194.325 100.640 196.385 ;
        RECT 102.800 194.325 102.940 197.065 ;
        RECT 104.110 195.765 104.390 195.880 ;
        RECT 104.640 195.765 104.780 197.745 ;
        RECT 107.400 197.385 107.540 199.105 ;
        RECT 108.780 197.725 108.920 213.385 ;
        RECT 109.640 211.685 109.900 212.005 ;
        RECT 109.180 207.605 109.440 207.925 ;
        RECT 109.240 206.565 109.380 207.605 ;
        RECT 109.180 206.245 109.440 206.565 ;
        RECT 109.180 203.525 109.440 203.845 ;
        RECT 109.240 201.125 109.380 203.525 ;
        RECT 109.700 202.825 109.840 211.685 ;
        RECT 112.460 208.120 112.600 216.105 ;
        RECT 113.780 215.485 114.040 215.745 ;
        RECT 113.380 215.425 114.040 215.485 ;
        RECT 113.380 215.345 113.980 215.425 ;
        RECT 113.380 213.025 113.520 215.345 ;
        RECT 117.450 215.230 117.730 215.600 ;
        RECT 122.980 215.425 123.240 215.745 ;
        RECT 123.900 215.425 124.160 215.745 ;
        RECT 117.520 214.045 117.660 215.230 ;
        RECT 121.600 214.405 121.860 214.725 ;
        RECT 114.240 213.725 114.500 214.045 ;
        RECT 117.460 213.725 117.720 214.045 ;
        RECT 120.210 213.870 120.490 214.240 ;
        RECT 120.220 213.725 120.480 213.870 ;
        RECT 112.860 212.705 113.120 213.025 ;
        RECT 113.320 212.880 113.580 213.025 ;
        RECT 112.920 210.840 113.060 212.705 ;
        RECT 113.310 212.510 113.590 212.880 ;
        RECT 112.850 210.470 113.130 210.840 ;
        RECT 110.090 207.750 110.370 208.120 ;
        RECT 112.390 207.750 112.670 208.120 ;
        RECT 110.160 202.825 110.300 207.750 ;
        RECT 112.920 205.885 113.060 210.470 ;
        RECT 113.380 210.045 113.520 212.510 ;
        RECT 114.300 212.005 114.440 213.725 ;
        RECT 114.240 211.685 114.500 212.005 ;
        RECT 117.520 210.985 117.660 213.725 ;
        RECT 120.220 213.045 120.480 213.365 ;
        RECT 120.280 211.325 120.420 213.045 ;
        RECT 121.140 212.705 121.400 213.025 ;
        RECT 121.200 211.325 121.340 212.705 ;
        RECT 118.380 211.005 118.640 211.325 ;
        RECT 120.220 211.005 120.480 211.325 ;
        RECT 121.140 211.005 121.400 211.325 ;
        RECT 117.460 210.665 117.720 210.985 ;
        RECT 114.230 210.045 114.510 210.160 ;
        RECT 113.380 209.905 114.510 210.045 ;
        RECT 114.230 209.790 114.510 209.905 ;
        RECT 115.610 207.750 115.890 208.120 ;
        RECT 116.540 207.945 116.800 208.265 ;
        RECT 115.620 207.605 115.880 207.750 ;
        RECT 116.600 207.585 116.740 207.945 ;
        RECT 117.460 207.605 117.720 207.925 ;
        RECT 116.540 207.265 116.800 207.585 ;
        RECT 112.860 205.565 113.120 205.885 ;
        RECT 113.310 205.710 113.590 206.080 ;
        RECT 116.600 205.965 116.740 207.265 ;
        RECT 114.760 205.885 116.740 205.965 ;
        RECT 114.240 205.795 114.500 205.885 ;
        RECT 114.760 205.825 116.800 205.885 ;
        RECT 114.760 205.795 114.900 205.825 ;
        RECT 111.020 205.225 111.280 205.545 ;
        RECT 109.640 202.505 109.900 202.825 ;
        RECT 110.100 202.505 110.360 202.825 ;
        RECT 109.700 201.320 109.840 202.505 ;
        RECT 109.180 200.805 109.440 201.125 ;
        RECT 109.630 200.950 109.910 201.320 ;
        RECT 108.720 197.405 108.980 197.725 ;
        RECT 107.340 197.065 107.600 197.385 ;
        RECT 105.040 196.385 105.300 196.705 ;
        RECT 105.500 196.385 105.760 196.705 ;
        RECT 106.420 196.560 106.680 196.705 ;
        RECT 105.100 195.880 105.240 196.385 ;
        RECT 104.110 195.625 104.780 195.765 ;
        RECT 104.110 195.510 104.390 195.625 ;
        RECT 105.030 195.510 105.310 195.880 ;
        RECT 103.660 194.685 103.920 195.005 ;
        RECT 104.580 194.685 104.840 195.005 ;
        RECT 100.440 194.005 100.700 194.325 ;
        RECT 102.740 194.005 103.000 194.325 ;
        RECT 102.280 193.665 102.540 193.985 ;
        RECT 103.200 193.665 103.460 193.985 ;
        RECT 102.340 192.285 102.480 193.665 ;
        RECT 102.280 191.965 102.540 192.285 ;
        RECT 103.260 191.945 103.400 193.665 ;
        RECT 99.520 191.625 99.780 191.945 ;
        RECT 103.200 191.625 103.460 191.945 ;
        RECT 99.060 191.285 99.320 191.605 ;
        RECT 99.580 189.225 99.720 191.625 ;
        RECT 101.360 190.945 101.620 191.265 ;
        RECT 101.420 189.510 101.560 190.945 ;
        RECT 103.720 190.245 103.860 194.685 ;
        RECT 104.120 193.840 104.380 193.985 ;
        RECT 104.110 193.470 104.390 193.840 ;
        RECT 104.640 192.285 104.780 194.685 ;
        RECT 104.580 191.965 104.840 192.285 ;
        RECT 105.100 191.945 105.240 195.510 ;
        RECT 105.560 194.665 105.700 196.385 ;
        RECT 106.410 196.190 106.690 196.560 ;
        RECT 109.240 195.005 109.380 200.805 ;
        RECT 109.630 200.270 109.910 200.640 ;
        RECT 109.700 198.405 109.840 200.270 ;
        RECT 111.080 199.960 111.220 205.225 ;
        RECT 113.380 204.865 113.520 205.710 ;
        RECT 114.240 205.655 114.900 205.795 ;
        RECT 114.240 205.565 114.500 205.655 ;
        RECT 116.540 205.565 116.800 205.825 ;
        RECT 113.770 205.030 114.050 205.400 ;
        RECT 113.320 204.545 113.580 204.865 ;
        RECT 113.840 203.505 113.980 205.030 ;
        RECT 114.300 204.040 114.440 205.565 ;
        RECT 115.620 205.455 115.880 205.545 ;
        RECT 115.620 205.315 116.280 205.455 ;
        RECT 115.620 205.225 115.880 205.315 ;
        RECT 114.230 203.670 114.510 204.040 ;
        RECT 113.780 203.360 114.040 203.505 ;
        RECT 111.480 202.845 111.740 203.165 ;
        RECT 113.770 202.990 114.050 203.360 ;
        RECT 110.560 199.445 110.820 199.765 ;
        RECT 111.010 199.590 111.290 199.960 ;
        RECT 109.640 198.085 109.900 198.405 ;
        RECT 109.640 197.405 109.900 197.725 ;
        RECT 105.960 194.685 106.220 195.005 ;
        RECT 109.180 194.685 109.440 195.005 ;
        RECT 105.500 194.345 105.760 194.665 ;
        RECT 105.040 191.625 105.300 191.945 ;
        RECT 103.660 189.925 103.920 190.245 ;
        RECT 106.020 189.510 106.160 194.685 ;
        RECT 109.700 194.665 109.840 197.405 ;
        RECT 110.620 197.385 110.760 199.445 ;
        RECT 111.540 199.425 111.680 202.845 ;
        RECT 112.860 202.505 113.120 202.825 ;
        RECT 114.240 202.505 114.500 202.825 ;
        RECT 114.700 202.680 114.960 202.825 ;
        RECT 112.920 199.960 113.060 202.505 ;
        RECT 114.300 201.320 114.440 202.505 ;
        RECT 114.690 202.310 114.970 202.680 ;
        RECT 115.620 202.165 115.880 202.485 ;
        RECT 114.230 200.950 114.510 201.320 ;
        RECT 115.680 200.105 115.820 202.165 ;
        RECT 116.140 200.105 116.280 205.315 ;
        RECT 117.000 205.225 117.260 205.545 ;
        RECT 117.060 203.845 117.200 205.225 ;
        RECT 117.520 205.205 117.660 207.605 ;
        RECT 117.460 204.885 117.720 205.205 ;
        RECT 118.440 203.845 118.580 211.005 ;
        RECT 120.680 210.665 120.940 210.985 ;
        RECT 119.300 209.985 119.560 210.305 ;
        RECT 119.760 209.985 120.020 210.305 ;
        RECT 118.830 208.430 119.110 208.800 ;
        RECT 118.900 208.265 119.040 208.430 ;
        RECT 118.840 207.945 119.100 208.265 ;
        RECT 119.360 207.585 119.500 209.985 ;
        RECT 119.300 207.265 119.560 207.585 ;
        RECT 119.360 205.205 119.500 207.265 ;
        RECT 119.820 206.565 119.960 209.985 ;
        RECT 120.220 207.265 120.480 207.585 ;
        RECT 119.760 206.245 120.020 206.565 ;
        RECT 119.300 204.885 119.560 205.205 ;
        RECT 117.000 203.525 117.260 203.845 ;
        RECT 118.380 203.525 118.640 203.845 ;
        RECT 116.540 202.505 116.800 202.825 ;
        RECT 116.600 200.445 116.740 202.505 ;
        RECT 117.060 202.485 117.200 203.525 ;
        RECT 117.000 202.165 117.260 202.485 ;
        RECT 118.440 200.445 118.580 203.525 ;
        RECT 118.840 202.165 119.100 202.485 ;
        RECT 116.540 200.125 116.800 200.445 ;
        RECT 118.380 200.125 118.640 200.445 ;
        RECT 112.850 199.590 113.130 199.960 ;
        RECT 115.620 199.785 115.880 200.105 ;
        RECT 116.080 199.785 116.340 200.105 ;
        RECT 111.480 199.105 111.740 199.425 ;
        RECT 110.560 197.065 110.820 197.385 ;
        RECT 111.020 197.065 111.280 197.385 ;
        RECT 110.550 195.510 110.830 195.880 ;
        RECT 111.080 195.685 111.220 197.065 ;
        RECT 112.400 196.725 112.660 197.045 ;
        RECT 111.940 196.385 112.200 196.705 ;
        RECT 110.620 195.005 110.760 195.510 ;
        RECT 111.020 195.365 111.280 195.685 ;
        RECT 110.560 194.915 110.820 195.005 ;
        RECT 110.160 194.775 110.820 194.915 ;
        RECT 109.640 194.345 109.900 194.665 ;
        RECT 110.160 192.965 110.300 194.775 ;
        RECT 110.560 194.685 110.820 194.775 ;
        RECT 111.480 194.685 111.740 195.005 ;
        RECT 112.000 194.915 112.140 196.385 ;
        RECT 112.460 195.685 112.600 196.725 ;
        RECT 113.780 196.385 114.040 196.705 ;
        RECT 112.400 195.365 112.660 195.685 ;
        RECT 113.840 195.005 113.980 196.385 ;
        RECT 115.680 195.685 115.820 199.785 ;
        RECT 115.620 195.365 115.880 195.685 ;
        RECT 116.540 195.025 116.800 195.345 ;
        RECT 112.400 194.915 112.660 195.005 ;
        RECT 112.000 194.775 112.660 194.915 ;
        RECT 112.400 194.685 112.660 194.775 ;
        RECT 113.780 194.685 114.040 195.005 ;
        RECT 115.620 194.685 115.880 195.005 ;
        RECT 111.540 193.985 111.680 194.685 ;
        RECT 111.480 193.665 111.740 193.985 ;
        RECT 112.460 193.840 112.600 194.685 ;
        RECT 115.680 194.520 115.820 194.685 ;
        RECT 115.610 194.150 115.890 194.520 ;
        RECT 112.390 193.470 112.670 193.840 ;
        RECT 110.100 192.645 110.360 192.965 ;
        RECT 110.560 192.645 110.820 192.965 ;
        RECT 101.420 189.370 106.160 189.510 ;
        RECT 99.520 188.905 99.780 189.225 ;
        RECT 101.420 187.715 101.560 189.370 ;
        RECT 106.020 187.715 106.160 189.370 ;
        RECT 110.620 188.810 110.760 192.645 ;
        RECT 116.600 192.625 116.740 195.025 ;
        RECT 118.900 194.665 119.040 202.165 ;
        RECT 119.360 194.665 119.500 204.885 ;
        RECT 119.820 204.865 119.960 206.245 ;
        RECT 120.280 206.225 120.420 207.265 ;
        RECT 120.740 206.565 120.880 210.665 ;
        RECT 121.660 208.685 121.800 214.405 ;
        RECT 122.060 213.725 122.320 214.045 ;
        RECT 121.200 208.545 121.800 208.685 ;
        RECT 120.680 206.245 120.940 206.565 ;
        RECT 120.220 205.905 120.480 206.225 ;
        RECT 121.200 204.865 121.340 208.545 ;
        RECT 121.600 207.605 121.860 207.925 ;
        RECT 121.660 206.225 121.800 207.605 ;
        RECT 121.600 205.905 121.860 206.225 ;
        RECT 122.120 205.885 122.260 213.725 ;
        RECT 123.040 213.365 123.180 215.425 ;
        RECT 123.960 213.365 124.100 215.425 ;
        RECT 122.980 213.045 123.240 213.365 ;
        RECT 123.900 213.045 124.160 213.365 ;
        RECT 122.520 211.345 122.780 211.665 ;
        RECT 122.060 205.565 122.320 205.885 ;
        RECT 119.760 204.545 120.020 204.865 ;
        RECT 121.140 204.720 121.400 204.865 ;
        RECT 121.130 204.350 121.410 204.720 ;
        RECT 122.060 202.845 122.320 203.165 ;
        RECT 122.120 201.125 122.260 202.845 ;
        RECT 122.060 200.805 122.320 201.125 ;
        RECT 121.140 200.465 121.400 200.785 ;
        RECT 121.200 200.105 121.340 200.465 ;
        RECT 121.140 199.785 121.400 200.105 ;
        RECT 119.760 196.725 120.020 197.045 ;
        RECT 119.820 195.005 119.960 196.725 ;
        RECT 119.760 194.915 120.020 195.005 ;
        RECT 119.760 194.775 120.420 194.915 ;
        RECT 119.760 194.685 120.020 194.775 ;
        RECT 118.380 194.345 118.640 194.665 ;
        RECT 118.840 194.345 119.100 194.665 ;
        RECT 119.300 194.345 119.560 194.665 ;
        RECT 117.920 193.665 118.180 193.985 ;
        RECT 117.980 193.160 118.120 193.665 ;
        RECT 117.910 192.790 118.190 193.160 ;
        RECT 118.440 192.965 118.580 194.345 ;
        RECT 119.360 193.895 119.500 194.345 ;
        RECT 118.900 193.755 119.500 193.895 ;
        RECT 118.380 192.645 118.640 192.965 ;
        RECT 116.540 192.305 116.800 192.625 ;
        RECT 115.160 191.285 115.420 191.605 ;
        RECT 113.780 190.945 114.040 191.265 ;
        RECT 113.840 189.565 113.980 190.945 ;
        RECT 113.780 189.245 114.040 189.565 ;
        RECT 115.220 188.810 115.360 191.285 ;
        RECT 110.620 188.670 115.360 188.810 ;
        RECT 110.620 187.840 110.760 188.670 ;
        RECT 96.750 187.160 97.030 187.715 ;
        RECT 92.150 187.020 97.030 187.160 ;
        RECT 92.150 185.715 92.430 187.020 ;
        RECT 96.750 186.290 97.030 187.020 ;
        RECT 96.690 185.890 97.030 186.290 ;
        RECT 96.750 185.715 97.030 185.890 ;
        RECT 101.350 185.715 101.630 187.715 ;
        RECT 105.950 186.690 106.230 187.715 ;
        RECT 110.540 187.440 110.840 187.840 ;
        RECT 115.220 187.715 115.360 188.670 ;
        RECT 118.900 188.155 119.040 193.755 ;
        RECT 119.760 192.645 120.020 192.965 ;
        RECT 119.300 191.965 119.560 192.285 ;
        RECT 119.360 189.905 119.500 191.965 ;
        RECT 119.300 189.585 119.560 189.905 ;
        RECT 119.820 188.660 119.960 192.645 ;
        RECT 120.280 192.285 120.420 194.775 ;
        RECT 121.200 193.160 121.340 199.785 ;
        RECT 122.120 195.345 122.260 200.805 ;
        RECT 122.580 197.725 122.720 211.345 ;
        RECT 123.040 203.360 123.180 213.045 ;
        RECT 123.440 205.795 123.700 205.885 ;
        RECT 123.960 205.795 124.100 213.045 ;
        RECT 124.880 212.005 125.020 216.445 ;
        RECT 127.640 216.085 127.780 216.445 ;
        RECT 125.740 215.765 126.000 216.085 ;
        RECT 127.580 215.765 127.840 216.085 ;
        RECT 125.280 212.705 125.540 213.025 ;
        RECT 124.820 211.685 125.080 212.005 ;
        RECT 125.340 211.665 125.480 212.705 ;
        RECT 125.280 211.345 125.540 211.665 ;
        RECT 125.800 209.285 125.940 215.765 ;
        RECT 128.040 215.425 128.300 215.745 ;
        RECT 127.580 213.725 127.840 214.045 ;
        RECT 127.120 213.385 127.380 213.705 ;
        RECT 125.740 208.965 126.000 209.285 ;
        RECT 127.180 208.945 127.320 213.385 ;
        RECT 127.640 210.985 127.780 213.725 ;
        RECT 128.100 213.705 128.240 215.425 ;
        RECT 128.040 213.385 128.300 213.705 ;
        RECT 127.580 210.665 127.840 210.985 ;
        RECT 127.570 209.790 127.850 210.160 ;
        RECT 127.120 208.625 127.380 208.945 ;
        RECT 127.120 207.265 127.380 207.585 ;
        RECT 126.200 205.905 126.460 206.225 ;
        RECT 123.440 205.655 124.100 205.795 ;
        RECT 123.440 205.565 123.700 205.655 ;
        RECT 125.280 205.565 125.540 205.885 ;
        RECT 122.970 202.990 123.250 203.360 ;
        RECT 123.500 200.445 123.640 205.565 ;
        RECT 124.360 204.545 124.620 204.865 ;
        RECT 124.420 202.145 124.560 204.545 ;
        RECT 125.340 203.360 125.480 205.565 ;
        RECT 125.270 202.990 125.550 203.360 ;
        RECT 124.880 202.485 125.940 202.565 ;
        RECT 124.880 202.425 126.000 202.485 ;
        RECT 124.360 201.825 124.620 202.145 ;
        RECT 124.880 201.125 125.020 202.425 ;
        RECT 125.740 202.165 126.000 202.425 ;
        RECT 124.820 200.805 125.080 201.125 ;
        RECT 123.440 200.125 123.700 200.445 ;
        RECT 123.500 199.425 123.640 200.125 ;
        RECT 126.260 199.765 126.400 205.905 ;
        RECT 126.660 201.825 126.920 202.145 ;
        RECT 126.200 199.445 126.460 199.765 ;
        RECT 123.440 199.105 123.700 199.425 ;
        RECT 123.500 198.065 123.640 199.105 ;
        RECT 123.440 197.745 123.700 198.065 ;
        RECT 122.520 197.405 122.780 197.725 ;
        RECT 126.200 197.065 126.460 197.385 ;
        RECT 123.900 196.725 124.160 197.045 ;
        RECT 122.060 195.025 122.320 195.345 ;
        RECT 123.960 194.665 124.100 196.725 ;
        RECT 124.360 196.385 124.620 196.705 ;
        RECT 123.900 194.345 124.160 194.665 ;
        RECT 122.970 193.470 123.250 193.840 ;
        RECT 121.130 192.790 121.410 193.160 ;
        RECT 120.220 191.965 120.480 192.285 ;
        RECT 121.200 191.605 121.340 192.790 ;
        RECT 123.040 191.945 123.180 193.470 ;
        RECT 122.980 191.625 123.240 191.945 ;
        RECT 121.140 191.285 121.400 191.605 ;
        RECT 121.200 189.225 121.340 191.285 ;
        RECT 121.140 188.905 121.400 189.225 ;
        RECT 124.420 188.660 124.560 196.385 ;
        RECT 126.260 195.685 126.400 197.065 ;
        RECT 126.200 195.365 126.460 195.685 ;
        RECT 126.720 195.005 126.860 201.825 ;
        RECT 127.180 196.705 127.320 207.265 ;
        RECT 127.640 205.885 127.780 209.790 ;
        RECT 128.560 206.225 128.700 216.445 ;
        RECT 131.720 213.725 131.980 214.045 ;
        RECT 130.340 213.385 130.600 213.705 ;
        RECT 128.960 211.345 129.220 211.665 ;
        RECT 129.020 208.120 129.160 211.345 ;
        RECT 130.400 210.305 130.540 213.385 ;
        RECT 130.340 209.985 130.600 210.305 ;
        RECT 129.880 208.965 130.140 209.285 ;
        RECT 129.420 208.625 129.680 208.945 ;
        RECT 128.950 207.750 129.230 208.120 ;
        RECT 128.960 207.605 129.220 207.750 ;
        RECT 129.480 206.565 129.620 208.625 ;
        RECT 129.940 206.565 130.080 208.965 ;
        RECT 130.400 208.605 130.540 209.985 ;
        RECT 130.340 208.285 130.600 208.605 ;
        RECT 129.420 206.245 129.680 206.565 ;
        RECT 129.880 206.245 130.140 206.565 ;
        RECT 128.500 205.905 128.760 206.225 ;
        RECT 127.580 205.565 127.840 205.885 ;
        RECT 128.560 205.545 128.700 205.905 ;
        RECT 129.940 205.885 130.080 206.245 ;
        RECT 128.960 205.565 129.220 205.885 ;
        RECT 129.880 205.565 130.140 205.885 ;
        RECT 130.340 205.565 130.600 205.885 ;
        RECT 131.260 205.565 131.520 205.885 ;
        RECT 128.500 205.225 128.760 205.545 ;
        RECT 128.560 203.505 128.700 205.225 ;
        RECT 128.500 203.185 128.760 203.505 ;
        RECT 128.500 202.505 128.760 202.825 ;
        RECT 128.560 200.640 128.700 202.505 ;
        RECT 127.580 200.125 127.840 200.445 ;
        RECT 128.490 200.270 128.770 200.640 ;
        RECT 129.020 200.445 129.160 205.565 ;
        RECT 129.870 202.990 130.150 203.360 ;
        RECT 129.940 202.825 130.080 202.990 ;
        RECT 129.880 202.505 130.140 202.825 ;
        RECT 129.420 201.825 129.680 202.145 ;
        RECT 129.480 200.785 129.620 201.825 ;
        RECT 129.940 200.785 130.080 202.505 ;
        RECT 129.420 200.465 129.680 200.785 ;
        RECT 129.880 200.465 130.140 200.785 ;
        RECT 128.960 200.125 129.220 200.445 ;
        RECT 127.640 198.405 127.780 200.125 ;
        RECT 128.490 199.590 128.770 199.960 ;
        RECT 128.040 199.105 128.300 199.425 ;
        RECT 127.580 198.085 127.840 198.405 ;
        RECT 128.100 197.385 128.240 199.105 ;
        RECT 128.040 197.065 128.300 197.385 ;
        RECT 127.120 196.385 127.380 196.705 ;
        RECT 128.040 196.385 128.300 196.705 ;
        RECT 128.100 195.880 128.240 196.385 ;
        RECT 128.030 195.510 128.310 195.880 ;
        RECT 126.660 194.685 126.920 195.005 ;
        RECT 125.280 192.305 125.540 192.625 ;
        RECT 125.740 192.305 126.000 192.625 ;
        RECT 125.340 190.245 125.480 192.305 ;
        RECT 125.800 191.265 125.940 192.305 ;
        RECT 128.560 191.945 128.700 199.590 ;
        RECT 129.480 197.385 129.620 200.465 ;
        RECT 129.420 197.065 129.680 197.385 ;
        RECT 128.950 195.510 129.230 195.880 ;
        RECT 128.960 195.365 129.220 195.510 ;
        RECT 130.400 194.325 130.540 205.565 ;
        RECT 130.800 201.825 131.060 202.145 ;
        RECT 130.860 201.125 131.000 201.825 ;
        RECT 130.800 200.805 131.060 201.125 ;
        RECT 131.320 195.005 131.460 205.565 ;
        RECT 131.780 205.400 131.920 213.725 ;
        RECT 133.100 213.045 133.360 213.365 ;
        RECT 133.160 212.005 133.300 213.045 ;
        RECT 132.640 211.685 132.900 212.005 ;
        RECT 133.100 211.685 133.360 212.005 ;
        RECT 132.700 207.585 132.840 211.685 ;
        RECT 133.620 208.605 133.760 218.825 ;
        RECT 134.470 218.265 134.750 223.050 ;
        RECT 146.400 222.750 146.700 222.900 ;
        RECT 146.400 222.500 146.710 222.750 ;
        RECT 143.220 219.505 143.480 219.825 ;
        RECT 134.540 216.765 134.680 218.265 ;
        RECT 140.920 218.145 141.180 218.465 ;
        RECT 139.530 217.270 139.810 217.640 ;
        RECT 134.480 216.445 134.740 216.765 ;
        RECT 134.020 216.105 134.280 216.425 ;
        RECT 134.080 213.365 134.220 216.105 ;
        RECT 134.480 215.765 134.740 216.085 ;
        RECT 135.390 215.910 135.670 216.280 ;
        RECT 136.780 216.105 137.040 216.425 ;
        RECT 139.080 216.105 139.340 216.425 ;
        RECT 134.020 213.045 134.280 213.365 ;
        RECT 134.540 210.305 134.680 215.765 ;
        RECT 135.460 211.325 135.600 215.910 ;
        RECT 135.860 212.705 136.120 213.025 ;
        RECT 135.400 211.005 135.660 211.325 ;
        RECT 135.920 210.985 136.060 212.705 ;
        RECT 136.840 212.200 136.980 216.105 ;
        RECT 138.620 215.425 138.880 215.745 ;
        RECT 138.160 213.045 138.420 213.365 ;
        RECT 136.770 211.830 137.050 212.200 ;
        RECT 135.860 210.665 136.120 210.985 ;
        RECT 134.480 209.985 134.740 210.305 ;
        RECT 133.560 208.285 133.820 208.605 ;
        RECT 134.020 207.605 134.280 207.925 ;
        RECT 132.640 207.265 132.900 207.585 ;
        RECT 131.710 205.030 131.990 205.400 ;
        RECT 133.560 205.225 133.820 205.545 ;
        RECT 132.180 204.885 132.440 205.205 ;
        RECT 132.640 204.885 132.900 205.205 ;
        RECT 131.710 200.270 131.990 200.640 ;
        RECT 131.780 199.425 131.920 200.270 ;
        RECT 131.720 199.105 131.980 199.425 ;
        RECT 131.780 197.385 131.920 199.105 ;
        RECT 131.720 197.065 131.980 197.385 ;
        RECT 132.240 196.705 132.380 204.885 ;
        RECT 132.700 200.640 132.840 204.885 ;
        RECT 133.100 204.545 133.360 204.865 ;
        RECT 133.160 201.125 133.300 204.545 ;
        RECT 133.100 200.805 133.360 201.125 ;
        RECT 132.630 200.270 132.910 200.640 ;
        RECT 132.630 198.230 132.910 198.600 ;
        RECT 132.700 198.065 132.840 198.230 ;
        RECT 132.640 197.745 132.900 198.065 ;
        RECT 131.720 196.385 131.980 196.705 ;
        RECT 132.180 196.385 132.440 196.705 ;
        RECT 131.260 194.685 131.520 195.005 ;
        RECT 128.960 194.005 129.220 194.325 ;
        RECT 130.340 194.005 130.600 194.325 ;
        RECT 129.020 192.285 129.160 194.005 ;
        RECT 131.320 192.625 131.460 194.685 ;
        RECT 131.260 192.305 131.520 192.625 ;
        RECT 131.780 192.480 131.920 196.385 ;
        RECT 132.630 196.190 132.910 196.560 ;
        RECT 132.700 195.345 132.840 196.190 ;
        RECT 133.160 195.595 133.300 200.805 ;
        RECT 133.620 200.105 133.760 205.225 ;
        RECT 134.080 202.485 134.220 207.605 ;
        RECT 134.020 202.165 134.280 202.485 ;
        RECT 133.560 199.785 133.820 200.105 ;
        RECT 134.080 195.685 134.220 202.165 ;
        RECT 134.540 200.105 134.680 209.985 ;
        RECT 135.400 207.265 135.660 207.585 ;
        RECT 134.940 200.125 135.200 200.445 ;
        RECT 134.480 199.785 134.740 200.105 ;
        RECT 133.160 195.455 133.760 195.595 ;
        RECT 132.640 195.025 132.900 195.345 ;
        RECT 133.620 195.005 133.760 195.455 ;
        RECT 134.020 195.365 134.280 195.685 ;
        RECT 134.480 195.365 134.740 195.685 ;
        RECT 133.100 194.685 133.360 195.005 ;
        RECT 133.560 194.685 133.820 195.005 ;
        RECT 132.640 194.345 132.900 194.665 ;
        RECT 132.700 192.625 132.840 194.345 ;
        RECT 133.160 193.160 133.300 194.685 ;
        RECT 133.560 194.005 133.820 194.325 ;
        RECT 133.090 192.790 133.370 193.160 ;
        RECT 128.960 191.965 129.220 192.285 ;
        RECT 131.710 192.110 131.990 192.480 ;
        RECT 132.640 192.305 132.900 192.625 ;
        RECT 128.040 191.625 128.300 191.945 ;
        RECT 128.500 191.625 128.760 191.945 ;
        RECT 125.740 190.945 126.000 191.265 ;
        RECT 128.100 191.120 128.240 191.625 ;
        RECT 133.160 191.265 133.300 192.790 ;
        RECT 128.030 190.750 128.310 191.120 ;
        RECT 129.420 190.945 129.680 191.265 ;
        RECT 133.100 190.945 133.360 191.265 ;
        RECT 129.480 190.465 129.620 190.945 ;
        RECT 129.020 190.325 129.620 190.465 ;
        RECT 125.280 189.925 125.540 190.245 ;
        RECT 119.820 188.520 124.560 188.660 ;
        RECT 118.840 187.835 119.100 188.155 ;
        RECT 119.820 187.715 119.960 188.520 ;
        RECT 124.420 187.715 124.560 188.520 ;
        RECT 129.020 187.715 129.160 190.325 ;
        RECT 133.620 188.960 133.760 194.005 ;
        RECT 134.080 192.285 134.220 195.365 ;
        RECT 134.540 194.520 134.680 195.365 ;
        RECT 135.000 195.005 135.140 200.125 ;
        RECT 134.940 194.685 135.200 195.005 ;
        RECT 134.470 194.150 134.750 194.520 ;
        RECT 134.020 191.965 134.280 192.285 ;
        RECT 134.540 191.945 134.680 194.150 ;
        RECT 135.460 191.945 135.600 207.265 ;
        RECT 137.240 206.245 137.500 206.565 ;
        RECT 137.300 200.445 137.440 206.245 ;
        RECT 136.320 200.125 136.580 200.445 ;
        RECT 137.240 200.125 137.500 200.445 ;
        RECT 136.380 199.845 136.520 200.125 ;
        RECT 136.380 199.705 137.440 199.845 ;
        RECT 137.300 199.425 137.440 199.705 ;
        RECT 136.780 199.105 137.040 199.425 ;
        RECT 137.240 199.105 137.500 199.425 ;
        RECT 136.320 196.725 136.580 197.045 ;
        RECT 134.480 191.625 134.740 191.945 ;
        RECT 135.400 191.625 135.660 191.945 ;
        RECT 135.860 191.625 136.120 191.945 ;
        RECT 135.920 189.565 136.060 191.625 ;
        RECT 136.380 189.760 136.520 196.725 ;
        RECT 136.840 195.005 136.980 199.105 ;
        RECT 138.220 197.125 138.360 213.045 ;
        RECT 138.680 212.005 138.820 215.425 ;
        RECT 139.140 213.025 139.280 216.105 ;
        RECT 139.080 212.705 139.340 213.025 ;
        RECT 138.620 211.685 138.880 212.005 ;
        RECT 139.140 211.520 139.280 212.705 ;
        RECT 139.070 211.150 139.350 211.520 ;
        RECT 139.600 208.265 139.740 217.270 ;
        RECT 140.980 216.765 141.120 218.145 ;
        RECT 143.280 217.445 143.420 219.505 ;
        RECT 144.130 219.310 144.410 219.680 ;
        RECT 141.840 217.125 142.100 217.445 ;
        RECT 143.220 217.125 143.480 217.445 ;
        RECT 141.900 216.960 142.040 217.125 ;
        RECT 140.920 216.445 141.180 216.765 ;
        RECT 141.830 216.590 142.110 216.960 ;
        RECT 144.200 216.765 144.340 219.310 ;
        RECT 145.060 219.165 145.320 219.485 ;
        RECT 144.140 216.445 144.400 216.765 ;
        RECT 140.000 216.105 140.260 216.425 ;
        RECT 140.060 214.725 140.200 216.105 ;
        RECT 140.000 214.405 140.260 214.725 ;
        RECT 144.590 214.550 144.870 214.920 ;
        RECT 143.670 213.870 143.950 214.240 ;
        RECT 140.920 213.385 141.180 213.705 ;
        RECT 142.760 213.385 143.020 213.705 ;
        RECT 140.000 212.705 140.260 213.025 ;
        RECT 140.060 211.665 140.200 212.705 ;
        RECT 140.980 212.200 141.120 213.385 ;
        RECT 140.910 212.085 141.190 212.200 ;
        RECT 140.520 211.945 141.190 212.085 ;
        RECT 140.000 211.345 140.260 211.665 ;
        RECT 140.000 210.665 140.260 210.985 ;
        RECT 139.540 207.945 139.800 208.265 ;
        RECT 139.080 207.265 139.340 207.585 ;
        RECT 139.140 205.885 139.280 207.265 ;
        RECT 139.080 205.565 139.340 205.885 ;
        RECT 140.060 202.565 140.200 210.665 ;
        RECT 139.600 202.425 140.200 202.565 ;
        RECT 138.620 201.825 138.880 202.145 ;
        RECT 137.760 196.985 138.360 197.125 ;
        RECT 137.240 196.385 137.500 196.705 ;
        RECT 136.780 194.685 137.040 195.005 ;
        RECT 137.300 191.800 137.440 196.385 ;
        RECT 137.760 192.625 137.900 196.985 ;
        RECT 138.160 196.385 138.420 196.705 ;
        RECT 138.220 193.840 138.360 196.385 ;
        RECT 138.150 193.470 138.430 193.840 ;
        RECT 138.160 192.645 138.420 192.965 ;
        RECT 137.700 192.305 137.960 192.625 ;
        RECT 137.230 191.430 137.510 191.800 ;
        RECT 138.220 189.760 138.360 192.645 ;
        RECT 135.860 189.245 136.120 189.565 ;
        RECT 136.310 189.390 136.590 189.760 ;
        RECT 138.150 189.390 138.430 189.760 ;
        RECT 138.680 189.165 138.820 201.825 ;
        RECT 139.080 200.125 139.340 200.445 ;
        RECT 139.140 199.425 139.280 200.125 ;
        RECT 139.600 199.765 139.740 202.425 ;
        RECT 140.000 201.825 140.260 202.145 ;
        RECT 139.540 199.445 139.800 199.765 ;
        RECT 139.080 199.105 139.340 199.425 ;
        RECT 139.600 198.405 139.740 199.445 ;
        RECT 139.540 198.085 139.800 198.405 ;
        RECT 139.540 197.065 139.800 197.385 ;
        RECT 139.080 196.385 139.340 196.705 ;
        RECT 139.140 192.480 139.280 196.385 ;
        RECT 139.070 192.110 139.350 192.480 ;
        RECT 138.220 189.025 138.820 189.165 ;
        RECT 138.220 188.960 138.360 189.025 ;
        RECT 133.620 188.820 138.360 188.960 ;
        RECT 133.620 187.715 133.760 188.820 ;
        RECT 138.220 187.715 138.360 188.820 ;
        RECT 139.600 188.495 139.740 197.065 ;
        RECT 140.060 196.560 140.200 201.825 ;
        RECT 139.990 196.190 140.270 196.560 ;
        RECT 140.520 194.665 140.660 211.945 ;
        RECT 140.910 211.830 141.190 211.945 ;
        RECT 141.840 210.160 142.100 210.305 ;
        RECT 141.830 209.790 142.110 210.160 ;
        RECT 141.840 207.265 142.100 207.585 ;
        RECT 141.900 206.080 142.040 207.265 ;
        RECT 142.820 206.760 142.960 213.385 ;
        RECT 143.740 213.025 143.880 213.870 ;
        RECT 143.680 212.705 143.940 213.025 ;
        RECT 144.660 211.325 144.800 214.550 ;
        RECT 144.600 211.005 144.860 211.325 ;
        RECT 144.590 209.110 144.870 209.480 ;
        RECT 143.680 208.800 143.940 208.945 ;
        RECT 143.670 208.430 143.950 208.800 ;
        RECT 144.660 208.265 144.800 209.110 ;
        RECT 144.600 207.945 144.860 208.265 ;
        RECT 142.750 206.390 143.030 206.760 ;
        RECT 140.920 205.565 141.180 205.885 ;
        RECT 141.830 205.710 142.110 206.080 ;
        RECT 144.140 205.565 144.400 205.885 ;
        RECT 140.980 202.000 141.120 205.565 ;
        RECT 141.840 204.545 142.100 204.865 ;
        RECT 141.900 203.360 142.040 204.545 ;
        RECT 141.830 202.990 142.110 203.360 ;
        RECT 140.910 201.630 141.190 202.000 ;
        RECT 143.220 201.825 143.480 202.145 ;
        RECT 143.680 202.000 143.940 202.145 ;
        RECT 141.380 200.805 141.640 201.125 ;
        RECT 140.920 200.125 141.180 200.445 ;
        RECT 140.980 199.280 141.120 200.125 ;
        RECT 140.910 198.910 141.190 199.280 ;
        RECT 140.920 194.685 141.180 195.005 ;
        RECT 140.460 194.345 140.720 194.665 ;
        RECT 140.980 192.965 141.120 194.685 ;
        RECT 140.920 192.645 141.180 192.965 ;
        RECT 141.440 192.365 141.580 200.805 ;
        RECT 143.280 200.445 143.420 201.825 ;
        RECT 143.670 201.630 143.950 202.000 ;
        RECT 143.220 200.125 143.480 200.445 ;
        RECT 141.840 199.105 142.100 199.425 ;
        RECT 143.680 199.105 143.940 199.425 ;
        RECT 141.900 197.920 142.040 199.105 ;
        RECT 141.830 197.550 142.110 197.920 ;
        RECT 143.740 197.725 143.880 199.105 ;
        RECT 143.680 197.405 143.940 197.725 ;
        RECT 142.760 197.240 143.020 197.385 ;
        RECT 142.750 196.870 143.030 197.240 ;
        RECT 141.840 196.385 142.100 196.705 ;
        RECT 143.680 196.560 143.940 196.705 ;
        RECT 141.900 193.840 142.040 196.385 ;
        RECT 143.670 196.190 143.950 196.560 ;
        RECT 143.210 195.510 143.490 195.880 ;
        RECT 143.280 195.005 143.420 195.510 ;
        RECT 143.220 194.685 143.480 195.005 ;
        RECT 143.680 194.345 143.940 194.665 ;
        RECT 141.830 193.470 142.110 193.840 ;
        RECT 142.760 193.665 143.020 193.985 ;
        RECT 140.980 192.225 141.580 192.365 ;
        RECT 140.980 191.945 141.120 192.225 ;
        RECT 140.920 191.625 141.180 191.945 ;
        RECT 142.300 191.625 142.560 191.945 ;
        RECT 141.840 190.945 142.100 191.265 ;
        RECT 141.900 189.905 142.040 190.945 ;
        RECT 141.840 189.585 142.100 189.905 ;
        RECT 139.540 188.175 139.800 188.495 ;
        RECT 142.360 188.155 142.500 191.625 ;
        RECT 142.300 187.835 142.560 188.155 ;
        RECT 142.820 187.715 142.960 193.665 ;
        RECT 143.740 190.245 143.880 194.345 ;
        RECT 143.680 189.925 143.940 190.245 ;
        RECT 144.200 188.885 144.340 205.565 ;
        RECT 145.120 202.825 145.260 219.165 ;
        RECT 145.510 217.950 145.790 218.320 ;
        RECT 146.430 218.265 146.710 222.500 ;
        RECT 149.590 219.540 149.890 219.640 ;
        RECT 150.600 219.540 150.900 219.690 ;
        RECT 149.590 219.390 150.900 219.540 ;
        RECT 149.590 219.240 149.890 219.390 ;
        RECT 150.600 219.290 150.900 219.390 ;
        RECT 145.580 217.445 145.720 217.950 ;
        RECT 145.520 217.125 145.780 217.445 ;
        RECT 145.970 215.230 146.250 215.600 ;
        RECT 146.040 213.025 146.180 215.230 ;
        RECT 146.500 214.045 146.640 218.265 ;
        RECT 149.590 218.240 149.890 218.290 ;
        RECT 151.000 218.240 151.300 218.390 ;
        RECT 149.590 218.090 151.300 218.240 ;
        RECT 149.590 217.890 149.890 218.090 ;
        RECT 151.000 217.990 151.300 218.090 ;
        RECT 149.590 216.890 149.890 216.940 ;
        RECT 151.350 216.890 151.650 217.040 ;
        RECT 149.590 216.740 151.650 216.890 ;
        RECT 149.590 216.540 149.890 216.740 ;
        RECT 151.350 216.640 151.650 216.740 ;
        RECT 149.590 215.490 149.890 215.590 ;
        RECT 151.650 215.490 151.950 215.640 ;
        RECT 149.590 215.340 151.950 215.490 ;
        RECT 149.590 215.190 149.890 215.340 ;
        RECT 151.650 215.240 151.950 215.340 ;
        RECT 149.590 214.140 149.890 214.190 ;
        RECT 151.950 214.140 152.250 214.290 ;
        RECT 146.440 213.725 146.700 214.045 ;
        RECT 149.590 213.990 152.250 214.140 ;
        RECT 149.590 213.790 149.890 213.990 ;
        RECT 151.950 213.890 152.250 213.990 ;
        RECT 145.510 212.510 145.790 212.880 ;
        RECT 145.980 212.705 146.240 213.025 ;
        RECT 149.590 212.740 149.890 212.790 ;
        RECT 152.250 212.740 152.550 212.890 ;
        RECT 149.590 212.590 152.550 212.740 ;
        RECT 145.580 212.005 145.720 212.510 ;
        RECT 149.590 212.390 149.890 212.590 ;
        RECT 152.250 212.490 152.550 212.590 ;
        RECT 145.520 211.685 145.780 212.005 ;
        RECT 145.510 211.150 145.790 211.520 ;
        RECT 149.590 211.440 149.890 211.490 ;
        RECT 152.550 211.440 152.850 211.590 ;
        RECT 149.590 211.290 152.850 211.440 ;
        RECT 145.580 209.285 145.720 211.150 ;
        RECT 149.590 211.090 149.890 211.290 ;
        RECT 152.550 211.190 152.850 211.290 ;
        RECT 149.590 210.090 149.890 210.140 ;
        RECT 152.850 210.090 153.150 210.240 ;
        RECT 149.590 209.940 153.150 210.090 ;
        RECT 149.590 209.740 149.890 209.940 ;
        RECT 152.850 209.840 153.150 209.940 ;
        RECT 145.520 208.965 145.780 209.285 ;
        RECT 149.590 208.690 149.890 208.790 ;
        RECT 153.150 208.690 153.450 208.840 ;
        RECT 149.590 208.540 153.450 208.690 ;
        RECT 149.590 208.390 149.890 208.540 ;
        RECT 153.150 208.440 153.450 208.540 ;
        RECT 145.510 207.070 145.790 207.440 ;
        RECT 149.590 207.340 149.890 207.390 ;
        RECT 153.450 207.340 153.750 207.490 ;
        RECT 149.590 207.190 153.750 207.340 ;
        RECT 145.580 206.565 145.720 207.070 ;
        RECT 149.590 206.990 149.890 207.190 ;
        RECT 153.450 207.090 153.750 207.190 ;
        RECT 145.520 206.245 145.780 206.565 ;
        RECT 149.590 206.040 149.890 206.090 ;
        RECT 153.750 206.040 154.050 206.190 ;
        RECT 149.590 205.890 154.050 206.040 ;
        RECT 149.590 205.690 149.890 205.890 ;
        RECT 153.750 205.790 154.050 205.890 ;
        RECT 145.510 204.350 145.790 204.720 ;
        RECT 149.590 204.640 149.890 204.740 ;
        RECT 154.050 204.640 154.350 204.790 ;
        RECT 149.590 204.490 154.350 204.640 ;
        RECT 145.580 203.845 145.720 204.350 ;
        RECT 149.590 204.340 149.890 204.490 ;
        RECT 154.050 204.390 154.350 204.490 ;
        RECT 145.520 203.525 145.780 203.845 ;
        RECT 149.590 203.290 149.890 203.390 ;
        RECT 154.350 203.290 154.650 203.440 ;
        RECT 149.590 203.140 154.650 203.290 ;
        RECT 149.590 202.990 149.890 203.140 ;
        RECT 154.350 203.040 154.650 203.140 ;
        RECT 145.060 202.505 145.320 202.825 ;
        RECT 149.590 201.890 149.890 201.990 ;
        RECT 154.650 201.890 154.950 202.040 ;
        RECT 149.590 201.740 154.950 201.890 ;
        RECT 149.590 201.590 149.890 201.740 ;
        RECT 154.650 201.640 154.950 201.740 ;
        RECT 145.510 200.270 145.790 200.640 ;
        RECT 149.590 200.590 149.890 200.690 ;
        RECT 154.950 200.590 155.250 200.740 ;
        RECT 149.590 200.440 155.250 200.590 ;
        RECT 149.590 200.290 149.890 200.440 ;
        RECT 154.950 200.340 155.250 200.440 ;
        RECT 145.580 199.765 145.720 200.270 ;
        RECT 145.520 199.445 145.780 199.765 ;
        RECT 145.510 198.910 145.790 199.280 ;
        RECT 149.590 199.240 149.890 199.290 ;
        RECT 155.250 199.240 155.550 199.390 ;
        RECT 149.590 199.090 155.550 199.240 ;
        RECT 145.580 198.405 145.720 198.910 ;
        RECT 149.590 198.890 149.890 199.090 ;
        RECT 155.250 198.990 155.550 199.090 ;
        RECT 145.520 198.085 145.780 198.405 ;
        RECT 149.590 197.890 149.890 197.940 ;
        RECT 155.550 197.890 155.850 198.040 ;
        RECT 149.590 197.740 155.850 197.890 ;
        RECT 149.590 197.540 149.890 197.740 ;
        RECT 155.550 197.640 155.850 197.740 ;
        RECT 149.590 196.440 149.890 196.540 ;
        RECT 155.850 196.440 156.150 196.590 ;
        RECT 149.590 196.290 156.150 196.440 ;
        RECT 149.590 196.140 149.890 196.290 ;
        RECT 155.850 196.190 156.150 196.290 ;
        RECT 145.520 195.365 145.780 195.685 ;
        RECT 145.580 195.200 145.720 195.365 ;
        RECT 144.590 194.830 144.870 195.200 ;
        RECT 145.510 194.830 145.790 195.200 ;
        RECT 149.640 195.090 149.940 195.190 ;
        RECT 156.150 195.090 156.450 195.240 ;
        RECT 149.625 194.940 156.450 195.090 ;
        RECT 144.600 194.685 144.860 194.830 ;
        RECT 149.640 194.790 149.940 194.940 ;
        RECT 156.150 194.840 156.450 194.940 ;
        RECT 149.590 193.790 149.890 193.890 ;
        RECT 156.450 193.790 156.750 193.940 ;
        RECT 149.590 193.640 156.750 193.790 ;
        RECT 149.590 193.490 149.890 193.640 ;
        RECT 156.450 193.540 156.750 193.640 ;
        RECT 149.590 192.340 149.890 192.440 ;
        RECT 156.750 192.340 157.050 192.490 ;
        RECT 149.590 192.190 157.050 192.340 ;
        RECT 149.590 192.040 149.890 192.190 ;
        RECT 156.750 192.090 157.050 192.190 ;
        RECT 147.360 191.285 147.620 191.605 ;
        RECT 144.140 188.565 144.400 188.885 ;
        RECT 147.420 187.715 147.560 191.285 ;
        RECT 149.590 190.990 149.890 191.140 ;
        RECT 157.050 190.990 157.350 191.140 ;
        RECT 149.590 190.840 157.350 190.990 ;
        RECT 149.590 190.740 149.890 190.840 ;
        RECT 157.050 190.740 157.350 190.840 ;
        RECT 149.540 189.590 149.840 189.740 ;
        RECT 157.350 189.590 157.650 189.740 ;
        RECT 149.540 189.440 157.650 189.590 ;
        RECT 149.540 189.340 149.840 189.440 ;
        RECT 157.350 189.340 157.650 189.440 ;
        RECT 105.940 186.290 106.240 186.690 ;
        RECT 105.950 185.715 106.230 186.290 ;
        RECT 110.550 185.715 110.830 187.440 ;
        RECT 115.150 185.715 115.430 187.715 ;
        RECT 119.750 187.490 120.030 187.715 ;
        RECT 119.740 187.090 120.040 187.490 ;
        RECT 119.750 185.715 120.030 187.090 ;
        RECT 124.350 185.715 124.630 187.715 ;
        RECT 128.950 186.690 129.230 187.715 ;
        RECT 133.550 187.140 133.830 187.715 ;
        RECT 133.540 186.740 133.840 187.140 ;
        RECT 128.940 186.290 129.240 186.690 ;
        RECT 128.950 185.715 129.230 186.290 ;
        RECT 133.550 185.715 133.830 186.740 ;
        RECT 138.150 185.715 138.430 187.715 ;
        RECT 142.750 186.690 143.030 187.715 ;
        RECT 142.740 186.290 143.040 186.690 ;
        RECT 145.840 186.290 146.140 186.690 ;
        RECT 142.750 185.715 143.030 186.290 ;
        RECT 41.590 185.390 41.740 185.715 ;
        RECT 41.490 184.990 41.790 185.390 ;
        RECT 14.640 182.340 15.490 182.840 ;
        RECT 7.290 181.945 7.590 182.085 ;
        RECT 7.290 181.795 8.340 181.945 ;
        RECT 7.290 181.685 7.590 181.795 ;
        RECT 8.190 181.645 8.340 181.795 ;
        RECT 8.115 181.245 8.415 181.645 ;
        RECT 16.490 180.940 17.340 182.740 ;
        RECT 25.465 182.145 25.765 182.255 ;
        RECT 18.315 181.995 25.765 182.145 ;
        RECT 18.315 181.845 18.465 181.995 ;
        RECT 25.465 181.855 25.765 181.995 ;
        RECT 18.265 181.445 18.565 181.845 ;
        RECT 20.965 181.145 21.265 181.295 ;
        RECT 25.465 181.145 25.765 181.205 ;
        RECT 20.965 180.995 25.765 181.145 ;
        RECT 20.965 180.895 21.265 180.995 ;
        RECT 7.290 180.745 7.590 180.885 ;
        RECT 25.465 180.805 25.765 180.995 ;
        RECT 10.865 180.745 11.165 180.795 ;
        RECT 7.290 180.595 11.165 180.745 ;
        RECT 7.290 180.485 7.590 180.595 ;
        RECT 10.865 180.395 11.165 180.595 ;
        RECT 6.915 179.615 7.215 179.755 ;
        RECT 6.915 179.495 8.440 179.615 ;
        RECT 16.490 179.590 17.340 180.090 ;
        RECT 25.090 179.565 25.390 179.675 ;
        RECT 6.915 179.465 8.465 179.495 ;
        RECT 6.915 179.355 7.215 179.465 ;
        RECT 8.165 179.095 8.465 179.465 ;
        RECT 18.340 179.415 25.390 179.565 ;
        RECT 18.340 179.195 18.490 179.415 ;
        RECT 25.090 179.275 25.390 179.415 ;
        RECT 6.540 178.815 6.840 178.955 ;
        RECT 6.540 178.665 11.515 178.815 ;
        RECT 6.540 178.555 6.840 178.665 ;
        RECT 11.365 178.515 11.515 178.665 ;
        RECT 14.065 178.515 14.365 178.915 ;
        RECT 18.265 178.795 18.565 179.195 ;
        RECT 24.715 179.020 25.015 179.130 ;
        RECT 20.390 178.870 25.015 179.020 ;
        RECT 20.390 178.590 20.540 178.870 ;
        RECT 24.715 178.730 25.015 178.870 ;
        RECT 6.915 178.165 7.215 178.305 ;
        RECT 10.815 178.165 11.115 178.295 ;
        RECT 6.915 178.015 11.115 178.165 ;
        RECT 11.365 178.115 11.665 178.515 ;
        RECT 6.915 177.905 7.215 178.015 ;
        RECT 10.815 177.895 11.115 178.015 ;
        RECT 6.540 177.565 6.840 177.705 ;
        RECT 14.140 177.565 14.290 178.515 ;
        RECT 15.065 178.465 20.540 178.590 ;
        RECT 15.015 178.440 20.540 178.465 ;
        RECT 15.015 178.065 15.315 178.440 ;
        RECT 20.965 178.415 21.265 178.515 ;
        RECT 25.090 178.415 25.390 178.475 ;
        RECT 20.965 178.265 25.390 178.415 ;
        RECT 17.665 177.845 17.965 178.245 ;
        RECT 20.965 178.115 21.265 178.265 ;
        RECT 25.090 178.075 25.390 178.265 ;
        RECT 26.940 178.390 27.240 178.490 ;
        RECT 32.615 178.390 32.915 178.440 ;
        RECT 35.640 178.390 35.940 178.490 ;
        RECT 26.940 178.190 35.940 178.390 ;
        RECT 26.940 178.090 27.240 178.190 ;
        RECT 32.615 178.040 32.915 178.190 ;
        RECT 35.640 178.090 35.940 178.190 ;
        RECT 6.540 177.415 14.290 177.565 ;
        RECT 17.740 177.665 17.890 177.845 ;
        RECT 24.715 177.665 25.015 177.725 ;
        RECT 17.740 177.515 25.015 177.665 ;
        RECT 6.540 177.305 6.840 177.415 ;
        RECT 14.640 176.890 15.490 177.390 ;
        RECT 24.715 177.325 25.015 177.515 ;
        RECT 24.340 176.905 24.640 177.015 ;
        RECT 18.315 176.755 24.640 176.905 ;
        RECT 6.170 176.505 6.470 176.645 ;
        RECT 6.170 176.355 8.340 176.505 ;
        RECT 18.315 176.405 18.465 176.755 ;
        RECT 24.340 176.615 24.640 176.755 ;
        RECT 6.170 176.245 6.470 176.355 ;
        RECT 8.190 176.205 8.340 176.355 ;
        RECT 8.115 175.805 8.415 176.205 ;
        RECT 5.790 175.655 6.090 175.795 ;
        RECT 11.365 175.755 11.665 176.155 ;
        RECT 15.015 175.830 15.315 176.205 ;
        RECT 18.265 176.005 18.565 176.405 ;
        RECT 23.965 176.330 24.265 176.440 ;
        RECT 18.740 176.180 24.265 176.330 ;
        RECT 18.740 175.830 18.890 176.180 ;
        RECT 23.965 176.040 24.265 176.180 ;
        RECT 35.640 176.040 35.940 176.140 ;
        RECT 15.015 175.805 18.890 175.830 ;
        RECT 11.365 175.655 11.515 175.755 ;
        RECT 5.790 175.505 11.515 175.655 ;
        RECT 5.790 175.395 6.090 175.505 ;
        RECT 14.065 175.355 14.365 175.755 ;
        RECT 15.065 175.680 18.890 175.805 ;
        RECT 20.965 175.705 21.265 175.855 ;
        RECT 34.370 175.840 35.940 176.040 ;
        RECT 24.340 175.705 24.640 175.765 ;
        RECT 35.640 175.740 35.940 175.840 ;
        RECT 20.965 175.555 24.640 175.705 ;
        RECT 20.965 175.455 21.265 175.555 ;
        RECT 6.170 175.140 6.470 175.280 ;
        RECT 10.865 175.140 11.165 175.355 ;
        RECT 6.170 174.990 11.165 175.140 ;
        RECT 6.170 174.880 6.470 174.990 ;
        RECT 10.865 174.955 11.165 174.990 ;
        RECT 5.790 174.620 6.090 174.760 ;
        RECT 14.115 174.620 14.265 175.355 ;
        RECT 17.715 175.055 18.015 175.455 ;
        RECT 24.340 175.365 24.640 175.555 ;
        RECT 23.965 175.055 24.265 175.115 ;
        RECT 17.715 174.905 24.265 175.055 ;
        RECT 23.965 174.715 24.265 174.905 ;
        RECT 5.790 174.470 14.265 174.620 ;
        RECT 5.790 174.360 6.090 174.470 ;
        RECT 16.490 174.140 17.340 174.640 ;
        RECT 23.590 174.125 23.890 174.235 ;
        RECT 36.340 174.190 37.140 180.440 ;
        RECT 37.540 180.090 39.390 182.740 ;
        RECT 50.790 182.640 50.940 185.715 ;
        RECT 55.390 183.090 55.540 185.715 ;
        RECT 64.590 184.040 64.740 185.715 ;
        RECT 73.790 184.490 73.940 185.715 ;
        RECT 82.990 184.940 83.140 185.715 ;
        RECT 82.940 184.540 83.240 184.940 ;
        RECT 105.290 184.690 105.590 184.840 ;
        RECT 108.740 184.690 109.040 184.840 ;
        RECT 105.290 184.540 109.040 184.690 ;
        RECT 73.740 184.090 74.040 184.490 ;
        RECT 105.290 184.440 105.590 184.540 ;
        RECT 108.740 184.440 109.040 184.540 ;
        RECT 64.540 183.640 64.840 184.040 ;
        RECT 104.840 183.440 105.140 183.590 ;
        RECT 107.940 183.440 108.240 183.590 ;
        RECT 104.840 183.290 108.240 183.440 ;
        RECT 104.840 183.190 105.140 183.290 ;
        RECT 107.940 183.190 108.240 183.290 ;
        RECT 55.290 182.690 55.590 183.090 ;
        RECT 103.390 182.990 103.690 183.140 ;
        RECT 108.390 182.990 108.690 183.140 ;
        RECT 103.390 182.840 108.690 182.990 ;
        RECT 103.390 182.740 103.690 182.840 ;
        RECT 108.390 182.740 108.690 182.840 ;
        RECT 50.740 182.240 51.040 182.640 ;
        RECT 76.140 180.940 77.990 182.740 ;
        RECT 115.240 180.940 117.090 185.540 ;
        RECT 73.220 180.530 73.520 180.580 ;
        RECT 84.970 180.530 85.320 180.580 ;
        RECT 38.640 178.365 38.940 178.540 ;
        RECT 38.165 178.215 38.940 178.365 ;
        RECT 5.420 173.980 5.720 174.120 ;
        RECT 8.165 173.980 8.465 174.055 ;
        RECT 5.420 173.830 8.465 173.980 ;
        RECT 5.420 173.720 5.720 173.830 ;
        RECT 8.165 173.655 8.465 173.830 ;
        RECT 18.340 173.975 23.890 174.125 ;
        RECT 38.165 174.140 38.315 178.215 ;
        RECT 38.640 178.140 38.940 178.215 ;
        RECT 38.640 175.740 38.940 176.140 ;
        RECT 38.715 174.690 38.865 175.740 ;
        RECT 39.890 175.440 40.190 180.440 ;
        RECT 41.140 180.040 44.240 180.440 ;
        RECT 41.490 177.540 41.790 180.040 ;
        RECT 43.540 177.540 43.890 180.040 ;
        RECT 40.540 177.140 40.840 177.240 ;
        RECT 41.990 177.140 42.290 177.240 ;
        RECT 40.540 176.940 42.290 177.140 ;
        RECT 40.540 176.840 40.840 176.940 ;
        RECT 41.990 176.840 42.290 176.940 ;
        RECT 43.090 177.140 43.390 177.240 ;
        RECT 44.540 177.140 44.840 177.240 ;
        RECT 43.090 176.940 44.840 177.140 ;
        RECT 43.090 176.840 43.390 176.940 ;
        RECT 44.540 176.840 44.840 176.940 ;
        RECT 45.190 175.440 45.490 180.440 ;
        RECT 70.270 180.230 85.320 180.530 ;
        RECT 70.270 179.880 70.620 180.230 ;
        RECT 73.220 180.180 73.520 180.230 ;
        RECT 84.970 180.130 85.320 180.230 ;
        RECT 59.920 178.580 102.920 179.080 ;
        RECT 67.420 178.530 67.720 178.580 ;
        RECT 83.870 178.180 84.170 178.280 ;
        RECT 83.870 177.980 103.670 178.180 ;
        RECT 83.870 177.880 84.170 177.980 ;
        RECT 78.770 177.580 79.070 177.680 ;
        RECT 81.640 177.580 81.940 177.690 ;
        RECT 78.770 177.380 103.670 177.580 ;
        RECT 78.770 177.280 79.070 177.380 ;
        RECT 81.640 177.290 81.940 177.380 ;
        RECT 71.020 176.930 71.320 177.080 ;
        RECT 72.270 176.930 72.570 177.080 ;
        RECT 71.020 176.780 72.570 176.930 ;
        RECT 71.020 176.680 71.320 176.780 ;
        RECT 72.270 176.680 72.570 176.780 ;
        RECT 71.420 176.430 71.720 176.580 ;
        RECT 72.770 176.430 73.070 176.580 ;
        RECT 73.570 176.430 78.170 176.830 ;
        RECT 71.420 176.280 73.070 176.430 ;
        RECT 71.420 176.180 71.720 176.280 ;
        RECT 72.770 176.180 73.070 176.280 ;
        RECT 86.570 176.080 102.920 176.580 ;
        RECT 73.920 175.480 83.220 175.880 ;
        RECT 85.870 175.730 86.170 175.780 ;
        RECT 98.140 175.730 98.440 175.790 ;
        RECT 99.490 175.730 99.790 175.790 ;
        RECT 103.170 175.730 103.470 175.780 ;
        RECT 85.870 175.430 103.470 175.730 ;
        RECT 85.870 175.380 86.170 175.430 ;
        RECT 98.140 175.390 98.440 175.430 ;
        RECT 99.490 175.390 99.790 175.430 ;
        RECT 103.170 175.380 103.470 175.430 ;
        RECT 40.990 174.690 41.290 174.840 ;
        RECT 42.790 174.690 43.090 174.840 ;
        RECT 38.715 174.540 43.090 174.690 ;
        RECT 40.990 174.440 41.290 174.540 ;
        RECT 42.790 174.440 43.090 174.540 ;
        RECT 74.345 174.480 97.170 175.030 ;
        RECT 42.290 174.140 42.590 174.290 ;
        RECT 44.090 174.140 44.390 174.290 ;
        RECT 38.165 173.990 44.390 174.140 ;
        RECT 18.340 173.755 18.490 173.975 ;
        RECT 23.590 173.835 23.890 173.975 ;
        RECT 42.290 173.890 42.590 173.990 ;
        RECT 44.090 173.890 44.390 173.990 ;
        RECT 51.820 174.230 52.120 174.330 ;
        RECT 70.970 174.230 71.270 174.330 ;
        RECT 87.240 174.230 87.540 174.340 ;
        RECT 51.820 174.030 87.540 174.230 ;
        RECT 51.820 173.930 52.120 174.030 ;
        RECT 70.970 173.930 71.270 174.030 ;
        RECT 87.240 173.940 87.540 174.030 ;
        RECT 108.690 174.015 108.990 174.110 ;
        RECT 125.195 174.015 125.495 184.815 ;
        RECT 142.240 184.640 145.040 185.490 ;
        RECT 145.890 184.840 146.040 186.290 ;
        RECT 147.350 185.715 147.630 187.715 ;
        RECT 148.040 185.990 148.340 186.390 ;
        RECT 147.440 184.840 147.590 185.715 ;
        RECT 148.140 184.840 148.290 185.990 ;
        RECT 145.790 184.440 146.090 184.840 ;
        RECT 147.440 184.440 147.740 184.840 ;
        RECT 148.040 184.440 148.340 184.840 ;
        RECT 150.090 184.290 150.390 184.440 ;
        RECT 143.445 184.140 150.390 184.290 ;
        RECT 143.445 183.915 143.595 184.140 ;
        RECT 150.090 184.040 150.390 184.140 ;
        RECT 143.345 183.515 143.645 183.915 ;
        RECT 144.145 183.815 144.495 183.965 ;
        RECT 145.795 183.815 146.095 183.965 ;
        RECT 144.145 183.665 149.495 183.815 ;
        RECT 144.145 183.515 144.495 183.665 ;
        RECT 145.795 183.565 146.095 183.665 ;
        RECT 142.045 183.365 142.345 183.415 ;
        RECT 146.295 183.365 146.595 183.515 ;
        RECT 142.045 183.215 146.595 183.365 ;
        RECT 142.045 183.015 142.345 183.215 ;
        RECT 146.295 183.115 146.595 183.215 ;
        RECT 143.695 182.965 143.995 183.065 ;
        RECT 146.745 182.965 147.045 183.065 ;
        RECT 143.695 182.815 147.045 182.965 ;
        RECT 143.695 182.665 143.995 182.815 ;
        RECT 146.745 182.665 147.045 182.815 ;
        RECT 142.145 181.600 142.445 181.750 ;
        RECT 147.145 181.600 147.445 181.800 ;
        RECT 142.145 181.450 147.445 181.600 ;
        RECT 142.145 181.350 142.445 181.450 ;
        RECT 147.145 181.400 147.445 181.450 ;
        RECT 147.990 181.215 148.290 181.290 ;
        RECT 143.395 181.065 149.495 181.215 ;
        RECT 143.395 180.865 143.545 181.065 ;
        RECT 147.990 180.890 148.290 181.065 ;
        RECT 143.295 180.465 143.595 180.865 ;
        RECT 144.145 180.665 144.495 180.865 ;
        RECT 145.795 180.665 146.095 180.865 ;
        RECT 144.145 180.515 146.095 180.665 ;
        RECT 144.145 180.415 144.495 180.515 ;
        RECT 145.795 180.465 146.095 180.515 ;
        RECT 143.345 180.215 143.645 180.315 ;
        RECT 145.395 180.215 145.695 180.315 ;
        RECT 143.345 180.065 145.695 180.215 ;
        RECT 143.345 179.915 143.645 180.065 ;
        RECT 145.395 179.915 145.695 180.065 ;
        RECT 144.545 179.615 144.895 179.665 ;
        RECT 148.895 179.615 149.245 179.665 ;
        RECT 144.545 179.265 149.245 179.615 ;
        RECT 144.545 179.215 144.895 179.265 ;
        RECT 148.895 179.215 149.245 179.265 ;
        RECT 142.145 178.565 142.445 178.965 ;
        RECT 143.845 178.915 144.145 179.065 ;
        RECT 148.045 178.915 148.345 179.065 ;
        RECT 143.845 178.765 148.345 178.915 ;
        RECT 143.845 178.665 144.145 178.765 ;
        RECT 148.045 178.665 148.345 178.765 ;
        RECT 142.195 178.415 142.345 178.565 ;
        RECT 148.445 178.415 148.745 178.515 ;
        RECT 142.195 178.265 148.745 178.415 ;
        RECT 148.445 178.115 148.745 178.265 ;
        RECT 143.245 177.915 143.560 178.095 ;
        RECT 143.245 177.865 143.645 177.915 ;
        RECT 147.545 177.865 147.845 177.915 ;
        RECT 143.245 177.715 147.845 177.865 ;
        RECT 143.245 177.665 143.560 177.715 ;
        RECT 143.495 177.115 143.795 177.515 ;
        RECT 144.745 177.165 145.045 177.565 ;
        RECT 147.545 177.515 147.845 177.715 ;
        RECT 142.545 176.115 142.845 176.165 ;
        RECT 143.545 176.115 143.695 177.115 ;
        RECT 142.545 175.915 143.695 176.115 ;
        RECT 143.895 176.115 144.245 176.215 ;
        RECT 144.795 176.115 144.995 177.165 ;
        RECT 143.895 175.915 144.995 176.115 ;
        RECT 142.545 175.765 142.845 175.915 ;
        RECT 143.895 175.815 144.245 175.915 ;
        RECT 143.495 175.265 143.795 175.415 ;
        RECT 145.845 175.265 146.145 175.415 ;
        RECT 143.495 175.115 146.145 175.265 ;
        RECT 143.495 175.015 143.795 175.115 ;
        RECT 145.845 175.015 146.145 175.115 ;
        RECT 142.095 174.615 142.395 174.765 ;
        RECT 147.145 174.615 147.445 174.765 ;
        RECT 142.095 174.415 147.445 174.615 ;
        RECT 142.095 174.365 142.395 174.415 ;
        RECT 147.145 174.365 147.445 174.415 ;
        RECT 144.195 174.165 144.545 174.215 ;
        RECT 148.895 174.165 149.245 174.215 ;
        RECT 79.740 173.880 80.040 173.890 ;
        RECT 79.720 173.780 80.040 173.880 ;
        RECT 5.040 173.375 5.340 173.515 ;
        RECT 5.040 173.225 11.515 173.375 ;
        RECT 5.040 173.115 5.340 173.225 ;
        RECT 11.365 173.075 11.515 173.225 ;
        RECT 14.065 173.075 14.365 173.475 ;
        RECT 18.265 173.355 18.565 173.755 ;
        RECT 23.215 173.580 23.515 173.690 ;
        RECT 20.390 173.430 23.515 173.580 ;
        RECT 78.370 173.580 80.040 173.780 ;
        RECT 108.690 173.815 128.795 174.015 ;
        RECT 108.690 173.710 108.990 173.815 ;
        RECT 125.195 173.765 125.495 173.815 ;
        RECT 78.370 173.430 78.570 173.580 ;
        RECT 79.720 173.490 80.040 173.580 ;
        RECT 102.490 173.530 105.140 173.540 ;
        RECT 79.720 173.480 80.020 173.490 ;
        RECT 20.390 173.150 20.540 173.430 ;
        RECT 23.215 173.290 23.515 173.430 ;
        RECT 5.420 172.725 5.720 172.865 ;
        RECT 10.815 172.725 11.115 172.855 ;
        RECT 5.420 172.575 11.115 172.725 ;
        RECT 11.365 172.675 11.665 173.075 ;
        RECT 5.420 172.465 5.720 172.575 ;
        RECT 10.815 172.455 11.115 172.575 ;
        RECT 5.040 172.125 5.340 172.265 ;
        RECT 14.140 172.125 14.290 173.075 ;
        RECT 15.065 173.025 20.540 173.150 ;
        RECT 40.640 173.190 40.940 173.390 ;
        RECT 44.440 173.215 44.740 173.390 ;
        RECT 15.015 173.000 20.540 173.025 ;
        RECT 15.015 172.625 15.315 173.000 ;
        RECT 20.965 172.975 21.265 173.075 ;
        RECT 40.640 173.040 41.665 173.190 ;
        RECT 23.590 172.975 23.890 173.035 ;
        RECT 20.965 172.825 23.890 172.975 ;
        RECT 17.665 172.405 17.965 172.805 ;
        RECT 20.965 172.675 21.265 172.825 ;
        RECT 23.590 172.635 23.890 172.825 ;
        RECT 26.505 172.940 26.805 173.020 ;
        RECT 33.240 172.940 33.540 173.040 ;
        RECT 35.690 172.940 35.990 173.040 ;
        RECT 26.505 172.740 35.990 172.940 ;
        RECT 26.505 172.620 26.805 172.740 ;
        RECT 33.240 172.640 33.540 172.740 ;
        RECT 35.690 172.640 35.990 172.740 ;
        RECT 37.240 172.640 37.540 173.040 ;
        RECT 40.640 172.990 40.940 173.040 ;
        RECT 5.040 171.975 14.290 172.125 ;
        RECT 17.740 172.225 17.890 172.405 ;
        RECT 23.215 172.225 23.515 172.285 ;
        RECT 17.740 172.075 23.515 172.225 ;
        RECT 5.040 171.865 5.340 171.975 ;
        RECT 14.640 171.440 15.490 171.940 ;
        RECT 23.215 171.885 23.515 172.075 ;
        RECT 22.840 171.465 23.140 171.575 ;
        RECT 18.315 171.315 23.140 171.465 ;
        RECT 4.670 171.065 4.970 171.205 ;
        RECT 4.670 170.915 8.340 171.065 ;
        RECT 18.315 170.965 18.465 171.315 ;
        RECT 22.840 171.175 23.140 171.315 ;
        RECT 4.670 170.805 4.970 170.915 ;
        RECT 8.190 170.765 8.340 170.915 ;
        RECT 8.115 170.365 8.415 170.765 ;
        RECT 4.290 170.215 4.590 170.355 ;
        RECT 11.365 170.315 11.665 170.715 ;
        RECT 15.015 170.390 15.315 170.765 ;
        RECT 18.265 170.565 18.565 170.965 ;
        RECT 22.465 170.890 22.765 171.000 ;
        RECT 18.740 170.740 22.765 170.890 ;
        RECT 37.340 170.790 37.540 172.640 ;
        RECT 18.740 170.390 18.890 170.740 ;
        RECT 22.465 170.600 22.765 170.740 ;
        RECT 15.015 170.365 18.890 170.390 ;
        RECT 11.365 170.215 11.515 170.315 ;
        RECT 4.290 170.065 11.515 170.215 ;
        RECT 4.290 169.955 4.590 170.065 ;
        RECT 14.065 169.915 14.365 170.315 ;
        RECT 15.065 170.240 18.890 170.365 ;
        RECT 20.965 170.265 21.265 170.415 ;
        RECT 37.290 170.390 37.590 170.790 ;
        RECT 22.840 170.265 23.140 170.325 ;
        RECT 20.965 170.115 23.140 170.265 ;
        RECT 20.965 170.015 21.265 170.115 ;
        RECT 4.670 169.700 4.970 169.840 ;
        RECT 10.865 169.700 11.165 169.915 ;
        RECT 4.670 169.550 11.165 169.700 ;
        RECT 4.670 169.440 4.970 169.550 ;
        RECT 10.865 169.515 11.165 169.550 ;
        RECT 4.290 169.180 4.590 169.320 ;
        RECT 14.115 169.180 14.265 169.915 ;
        RECT 17.715 169.615 18.015 170.015 ;
        RECT 22.840 169.925 23.140 170.115 ;
        RECT 39.940 169.890 40.240 172.790 ;
        RECT 41.515 172.240 41.665 173.040 ;
        RECT 43.740 173.065 44.740 173.215 ;
        RECT 43.740 172.240 43.890 173.065 ;
        RECT 44.440 172.990 44.740 173.065 ;
        RECT 41.490 171.840 41.790 172.240 ;
        RECT 43.640 171.840 43.940 172.240 ;
        RECT 40.490 171.040 40.790 171.440 ;
        RECT 40.540 170.240 40.690 171.040 ;
        RECT 41.540 170.240 41.740 171.840 ;
        RECT 43.690 170.240 43.890 171.840 ;
        RECT 44.540 171.040 44.840 171.440 ;
        RECT 44.640 170.240 44.790 171.040 ;
        RECT 40.490 169.840 40.790 170.240 ;
        RECT 41.490 169.840 41.790 170.240 ;
        RECT 43.640 169.840 43.940 170.240 ;
        RECT 44.540 169.840 44.840 170.240 ;
        RECT 45.240 169.890 45.540 172.790 ;
        RECT 61.320 172.730 71.320 173.130 ;
        RECT 78.320 173.030 78.620 173.430 ;
        RECT 86.570 173.040 105.140 173.530 ;
        RECT 86.570 173.030 102.920 173.040 ;
        RECT 74.345 172.240 97.190 172.790 ;
        RECT 71.020 171.630 78.170 172.030 ;
        RECT 66.670 171.330 66.970 171.430 ;
        RECT 72.270 171.330 72.570 171.430 ;
        RECT 66.670 171.130 72.570 171.330 ;
        RECT 66.670 171.030 66.970 171.130 ;
        RECT 72.270 171.030 72.570 171.130 ;
        RECT 48.270 170.880 48.570 170.980 ;
        RECT 48.270 170.680 68.820 170.880 ;
        RECT 48.270 170.580 48.570 170.680 ;
        RECT 43.040 169.690 43.340 169.790 ;
        RECT 46.890 169.690 47.190 169.740 ;
        RECT 22.465 169.615 22.765 169.675 ;
        RECT 17.715 169.465 22.765 169.615 ;
        RECT 22.465 169.275 22.765 169.465 ;
        RECT 43.040 169.490 47.190 169.690 ;
        RECT 43.040 169.390 43.340 169.490 ;
        RECT 46.890 169.340 47.190 169.490 ;
        RECT 4.290 169.030 14.265 169.180 ;
        RECT 4.290 168.920 4.590 169.030 ;
        RECT 16.490 168.740 17.340 169.240 ;
        RECT 22.090 168.685 22.390 168.795 ;
        RECT 3.920 168.540 4.220 168.680 ;
        RECT 8.165 168.540 8.465 168.615 ;
        RECT 3.920 168.390 8.465 168.540 ;
        RECT 3.920 168.280 4.220 168.390 ;
        RECT 8.165 168.215 8.465 168.390 ;
        RECT 18.340 168.535 22.390 168.685 ;
        RECT 18.340 168.315 18.490 168.535 ;
        RECT 22.090 168.395 22.390 168.535 ;
        RECT 40.940 168.540 41.240 168.640 ;
        RECT 42.490 168.540 42.790 168.640 ;
        RECT 44.090 168.540 44.390 168.640 ;
        RECT 40.940 168.340 44.390 168.540 ;
        RECT 3.540 167.935 3.840 168.075 ;
        RECT 3.540 167.785 11.515 167.935 ;
        RECT 3.540 167.675 3.840 167.785 ;
        RECT 11.365 167.635 11.515 167.785 ;
        RECT 14.065 167.635 14.365 168.035 ;
        RECT 18.265 167.915 18.565 168.315 ;
        RECT 21.715 168.140 22.015 168.250 ;
        RECT 40.940 168.240 41.240 168.340 ;
        RECT 42.490 168.240 42.790 168.340 ;
        RECT 44.090 168.240 44.390 168.340 ;
        RECT 51.020 168.280 51.220 170.680 ;
        RECT 68.420 170.580 68.820 170.680 ;
        RECT 70.370 170.680 70.670 170.780 ;
        RECT 86.470 170.680 86.770 170.830 ;
        RECT 70.370 170.530 86.770 170.680 ;
        RECT 67.820 170.480 68.220 170.530 ;
        RECT 54.120 170.280 68.220 170.480 ;
        RECT 70.370 170.380 70.670 170.530 ;
        RECT 86.470 170.430 86.770 170.530 ;
        RECT 54.120 170.080 54.420 170.280 ;
        RECT 67.820 170.230 68.220 170.280 ;
        RECT 61.820 169.630 83.220 170.030 ;
        RECT 92.420 169.830 92.720 170.230 ;
        RECT 93.720 170.080 94.020 170.230 ;
        RECT 103.170 170.080 103.470 170.230 ;
        RECT 93.720 169.930 103.470 170.080 ;
        RECT 93.720 169.830 94.020 169.930 ;
        RECT 103.170 169.830 103.470 169.930 ;
        RECT 92.495 169.480 92.645 169.830 ;
        RECT 54.470 169.330 92.645 169.480 ;
        RECT 98.870 169.330 99.170 169.430 ;
        RECT 101.820 169.330 102.120 169.430 ;
        RECT 54.470 169.080 62.770 169.330 ;
        RECT 98.870 169.290 103.670 169.330 ;
        RECT 103.890 169.290 104.190 169.440 ;
        RECT 54.470 168.830 54.870 169.080 ;
        RECT 64.770 169.030 65.070 169.180 ;
        RECT 98.870 169.140 104.190 169.290 ;
        RECT 98.870 169.130 103.670 169.140 ;
        RECT 67.220 169.030 67.520 169.130 ;
        RECT 64.770 168.980 67.520 169.030 ;
        RECT 86.220 168.980 86.520 169.080 ;
        RECT 88.320 168.980 88.620 169.080 ;
        RECT 98.870 169.030 99.170 169.130 ;
        RECT 101.820 169.030 102.120 169.130 ;
        RECT 103.890 169.040 104.190 169.140 ;
        RECT 51.520 168.430 54.870 168.830 ;
        RECT 55.270 168.530 61.620 168.930 ;
        RECT 64.770 168.880 88.620 168.980 ;
        RECT 64.770 168.780 65.070 168.880 ;
        RECT 67.220 168.780 88.620 168.880 ;
        RECT 67.220 168.730 67.520 168.780 ;
        RECT 86.220 168.680 86.520 168.780 ;
        RECT 88.320 168.680 88.620 168.780 ;
        RECT 94.370 168.880 94.670 169.030 ;
        RECT 104.890 168.890 105.140 173.040 ;
        RECT 108.240 169.565 108.540 169.660 ;
        RECT 125.195 169.565 125.495 173.165 ;
        RECT 128.595 171.615 128.795 173.815 ;
        RECT 144.195 173.815 149.245 174.165 ;
        RECT 144.195 173.765 144.545 173.815 ;
        RECT 148.895 173.765 149.245 173.815 ;
        RECT 145.845 173.515 146.145 173.665 ;
        RECT 147.995 173.515 148.295 173.665 ;
        RECT 145.845 173.365 148.295 173.515 ;
        RECT 145.845 173.265 146.145 173.365 ;
        RECT 147.995 173.265 148.295 173.365 ;
        RECT 143.645 173.115 143.945 173.265 ;
        RECT 146.695 173.115 146.995 173.215 ;
        RECT 143.645 172.965 146.995 173.115 ;
        RECT 143.645 172.865 143.945 172.965 ;
        RECT 146.695 172.815 146.995 172.965 ;
        RECT 142.645 172.215 142.995 172.315 ;
        RECT 145.845 172.215 146.145 172.315 ;
        RECT 142.645 172.015 146.145 172.215 ;
        RECT 142.645 171.865 142.995 172.015 ;
        RECT 145.845 171.915 146.145 172.015 ;
        RECT 139.445 171.615 139.745 171.715 ;
        RECT 142.385 171.615 142.685 171.725 ;
        RECT 128.595 171.415 142.685 171.615 ;
        RECT 139.445 171.315 139.745 171.415 ;
        RECT 142.385 171.325 142.685 171.415 ;
        RECT 142.925 171.615 143.225 171.725 ;
        RECT 144.895 171.615 145.195 171.715 ;
        RECT 142.925 171.415 145.195 171.615 ;
        RECT 142.925 171.325 143.225 171.415 ;
        RECT 144.895 171.315 145.195 171.415 ;
        RECT 148.295 171.315 148.595 171.715 ;
        RECT 142.145 171.065 142.445 171.165 ;
        RECT 147.545 171.065 147.845 171.215 ;
        RECT 142.145 170.915 149.495 171.065 ;
        RECT 142.145 170.765 142.445 170.915 ;
        RECT 147.545 170.815 147.845 170.915 ;
        RECT 141.345 170.615 141.645 170.715 ;
        RECT 144.445 170.615 144.745 170.715 ;
        RECT 141.345 170.415 144.745 170.615 ;
        RECT 141.345 170.315 141.645 170.415 ;
        RECT 144.445 170.315 144.745 170.415 ;
        RECT 143.145 170.115 143.445 170.215 ;
        RECT 145.295 170.115 145.595 170.265 ;
        RECT 143.145 169.965 145.595 170.115 ;
        RECT 143.145 169.815 143.445 169.965 ;
        RECT 145.295 169.865 145.595 169.965 ;
        RECT 142.385 169.565 142.685 169.665 ;
        RECT 108.240 169.365 142.685 169.565 ;
        RECT 108.240 169.260 108.540 169.365 ;
        RECT 94.370 168.740 104.365 168.880 ;
        RECT 94.370 168.730 104.440 168.740 ;
        RECT 94.370 168.630 94.670 168.730 ;
        RECT 85.670 168.530 85.970 168.630 ;
        RECT 86.720 168.530 87.020 168.630 ;
        RECT 87.770 168.530 88.070 168.630 ;
        RECT 88.820 168.530 89.120 168.630 ;
        RECT 89.870 168.530 90.170 168.630 ;
        RECT 20.390 167.990 22.015 168.140 ;
        RECT 20.390 167.710 20.540 167.990 ;
        RECT 21.715 167.850 22.015 167.990 ;
        RECT 41.990 168.040 42.290 168.140 ;
        RECT 48.870 168.130 57.020 168.280 ;
        RECT 62.420 168.130 64.320 168.530 ;
        RECT 85.670 168.330 90.170 168.530 ;
        RECT 85.670 168.230 85.970 168.330 ;
        RECT 86.720 168.230 87.020 168.330 ;
        RECT 87.770 168.230 88.070 168.330 ;
        RECT 88.820 168.230 89.120 168.330 ;
        RECT 89.870 168.230 90.170 168.330 ;
        RECT 93.070 168.430 93.370 168.580 ;
        RECT 93.070 168.280 103.865 168.430 ;
        RECT 104.140 168.340 104.440 168.730 ;
        RECT 93.070 168.180 93.370 168.280 ;
        RECT 46.565 168.040 57.020 168.130 ;
        RECT 41.990 167.980 57.020 168.040 ;
        RECT 41.990 167.840 46.790 167.980 ;
        RECT 48.870 167.880 57.020 167.980 ;
        RECT 41.990 167.740 42.290 167.840 ;
        RECT 3.920 167.285 4.220 167.425 ;
        RECT 10.815 167.285 11.115 167.415 ;
        RECT 3.920 167.135 11.115 167.285 ;
        RECT 11.365 167.235 11.665 167.635 ;
        RECT 3.920 167.025 4.220 167.135 ;
        RECT 10.815 167.015 11.115 167.135 ;
        RECT 3.540 166.685 3.840 166.825 ;
        RECT 14.140 166.685 14.290 167.635 ;
        RECT 15.065 167.585 20.540 167.710 ;
        RECT 15.015 167.560 20.540 167.585 ;
        RECT 15.015 167.185 15.315 167.560 ;
        RECT 20.965 167.535 21.265 167.635 ;
        RECT 22.090 167.535 22.390 167.595 ;
        RECT 20.965 167.385 22.390 167.535 ;
        RECT 17.665 166.965 17.965 167.365 ;
        RECT 20.965 167.235 21.265 167.385 ;
        RECT 22.090 167.195 22.390 167.385 ;
        RECT 46.890 167.580 47.190 167.690 ;
        RECT 51.970 167.580 60.070 167.680 ;
        RECT 63.570 167.580 66.820 167.980 ;
        RECT 73.220 167.930 73.520 168.080 ;
        RECT 100.420 167.930 100.720 168.080 ;
        RECT 67.220 167.730 67.520 167.880 ;
        RECT 68.920 167.730 69.220 167.880 ;
        RECT 70.520 167.730 70.820 167.880 ;
        RECT 67.220 167.580 70.820 167.730 ;
        RECT 73.220 167.780 100.720 167.930 ;
        RECT 103.715 167.965 103.865 168.280 ;
        RECT 104.140 167.965 104.440 168.090 ;
        RECT 103.715 167.815 104.440 167.965 ;
        RECT 73.220 167.680 73.520 167.780 ;
        RECT 100.420 167.680 100.720 167.780 ;
        RECT 104.140 167.690 104.440 167.815 ;
        RECT 46.890 167.430 60.070 167.580 ;
        RECT 67.220 167.480 67.520 167.580 ;
        RECT 68.920 167.480 69.220 167.580 ;
        RECT 70.520 167.480 70.820 167.580 ;
        RECT 104.890 167.490 107.990 168.890 ;
        RECT 108.240 168.340 108.540 168.740 ;
        RECT 108.590 167.690 108.890 168.090 ;
        RECT 46.890 167.290 47.190 167.430 ;
        RECT 51.970 167.280 60.070 167.430 ;
        RECT 62.420 167.230 65.320 167.380 ;
        RECT 95.270 167.230 95.570 167.380 ;
        RECT 3.540 166.535 14.290 166.685 ;
        RECT 17.740 166.785 17.890 166.965 ;
        RECT 21.715 166.785 22.015 166.845 ;
        RECT 17.740 166.635 22.015 166.785 ;
        RECT 48.420 166.730 57.920 167.130 ;
        RECT 58.320 166.730 62.170 167.130 ;
        RECT 62.420 167.080 95.595 167.230 ;
        RECT 62.420 166.980 65.320 167.080 ;
        RECT 95.270 166.980 95.570 167.080 ;
        RECT 3.540 166.425 3.840 166.535 ;
        RECT 14.640 165.990 15.490 166.490 ;
        RECT 21.715 166.445 22.015 166.635 ;
        RECT 57.520 166.480 57.920 166.730 ;
        RECT 64.270 166.530 64.570 166.680 ;
        RECT 67.220 166.530 67.520 166.680 ;
        RECT 57.520 166.080 62.770 166.480 ;
        RECT 64.270 166.380 67.520 166.530 ;
        RECT 64.270 166.280 64.570 166.380 ;
        RECT 67.220 166.280 67.520 166.380 ;
        RECT 72.520 166.630 72.820 166.680 ;
        RECT 98.870 166.630 99.170 166.730 ;
        RECT 72.520 166.430 99.170 166.630 ;
        RECT 72.520 166.280 72.820 166.430 ;
        RECT 98.870 166.330 99.170 166.430 ;
        RECT 39.640 164.190 41.340 165.990 ;
        RECT 66.890 164.190 68.590 165.990 ;
        RECT 105.240 163.640 105.540 164.040 ;
        RECT 77.465 161.340 77.765 161.740 ;
        RECT 77.915 161.640 78.215 162.040 ;
        RECT 78.365 161.940 78.665 162.340 ;
        RECT 78.815 162.240 79.115 162.640 ;
        RECT 79.265 162.540 79.565 162.940 ;
        RECT 79.715 162.840 80.015 163.240 ;
        RECT 32.640 160.245 34.340 160.290 ;
        RECT 20.205 159.780 37.550 160.245 ;
        RECT 10.290 158.840 10.590 158.890 ;
        RECT 10.290 158.790 10.665 158.840 ;
        RECT 19.940 158.790 20.940 159.235 ;
        RECT 21.500 158.895 22.500 159.780 ;
        RECT 32.640 159.740 34.340 159.780 ;
        RECT 27.045 159.505 27.920 159.610 ;
        RECT 41.395 159.505 42.270 159.565 ;
        RECT 27.045 159.350 42.270 159.505 ;
        RECT 27.920 159.345 42.270 159.350 ;
        RECT 10.290 158.590 20.940 158.790 ;
        RECT 23.195 158.810 31.935 158.870 ;
        RECT 23.195 158.610 31.940 158.810 ;
        RECT 10.290 158.540 10.665 158.590 ;
        RECT 10.290 158.490 10.590 158.540 ;
        RECT 19.940 158.235 20.940 158.590 ;
        RECT 26.965 158.275 27.965 158.330 ;
        RECT 3.290 157.890 3.590 157.990 ;
        RECT 26.860 157.890 28.110 158.275 ;
        RECT 31.680 157.935 31.940 158.610 ;
        RECT 38.420 158.420 38.680 158.700 ;
        RECT 39.380 158.420 39.640 158.700 ;
        RECT 40.340 158.420 40.600 158.700 ;
        RECT 38.420 158.160 40.600 158.420 ;
        RECT 3.290 157.690 28.110 157.890 ;
        RECT 3.290 157.590 3.590 157.690 ;
        RECT 20.670 156.990 23.590 157.460 ;
        RECT 26.860 157.400 28.110 157.690 ;
        RECT 26.965 157.330 27.965 157.400 ;
        RECT 32.870 157.390 33.130 157.820 ;
        RECT 34.210 157.390 34.470 157.830 ;
        RECT 36.285 157.390 37.285 157.930 ;
        RECT 38.420 157.825 38.680 158.160 ;
        RECT 39.380 157.825 39.640 158.160 ;
        RECT 40.340 157.825 40.600 158.160 ;
        RECT 38.860 157.390 39.120 157.670 ;
        RECT 39.820 157.390 40.080 157.670 ;
        RECT 32.870 157.360 40.080 157.390 ;
        RECT 40.995 157.360 41.155 159.345 ;
        RECT 41.395 159.305 42.270 159.345 ;
        RECT 43.905 159.250 44.780 159.510 ;
        RECT 32.870 157.200 41.155 157.360 ;
        RECT 32.870 157.130 40.080 157.200 ;
        RECT 5.240 154.570 5.590 154.790 ;
        RECT 20.670 154.570 21.125 156.990 ;
        RECT 25.280 156.630 25.540 157.060 ;
        RECT 27.330 156.630 27.590 157.010 ;
        RECT 32.870 156.945 33.130 157.130 ;
        RECT 34.210 156.955 34.470 157.130 ;
        RECT 36.285 156.930 37.285 157.130 ;
        RECT 38.860 156.795 39.120 157.130 ;
        RECT 39.820 156.795 40.080 157.130 ;
        RECT 44.135 156.630 44.635 159.250 ;
        RECT 55.285 159.240 56.160 159.500 ;
        RECT 61.185 159.240 62.060 159.500 ;
        RECT 70.045 159.240 70.920 159.500 ;
        RECT 25.280 156.380 44.635 156.630 ;
        RECT 21.410 155.240 22.410 156.240 ;
        RECT 25.280 156.185 25.540 156.380 ;
        RECT 27.330 156.135 27.590 156.380 ;
        RECT 23.515 155.155 23.775 156.030 ;
        RECT 29.480 155.850 29.740 156.190 ;
        RECT 35.400 155.850 35.660 156.190 ;
        RECT 29.480 155.610 35.660 155.850 ;
        RECT 29.480 155.315 29.740 155.610 ;
        RECT 35.400 155.315 35.660 155.610 ;
        RECT 23.585 154.980 23.735 155.155 ;
        RECT 29.945 154.980 37.000 155.165 ;
        RECT 41.380 155.085 41.640 155.960 ;
        RECT 44.135 155.240 44.635 156.380 ;
        RECT 55.485 155.240 55.985 159.240 ;
        RECT 61.435 155.240 61.935 159.240 ;
        RECT 70.235 155.240 70.735 159.240 ;
        RECT 23.585 154.965 39.865 154.980 ;
        RECT 23.585 154.780 30.185 154.965 ;
        RECT 36.755 154.780 39.865 154.965 ;
        RECT 24.935 154.710 25.810 154.780 ;
        RECT 29.120 154.710 30.185 154.780 ;
        RECT 21.665 154.570 22.665 154.695 ;
        RECT 31.755 154.570 32.630 154.675 ;
        RECT 35.080 154.570 35.955 154.675 ;
        RECT 38.860 154.665 39.865 154.780 ;
        RECT 41.435 154.570 41.585 155.085 ;
        RECT 43.885 154.980 44.760 155.240 ;
        RECT 55.235 154.980 56.110 155.240 ;
        RECT 61.135 154.980 62.010 155.240 ;
        RECT 70.035 154.980 70.910 155.240 ;
        RECT 5.240 154.305 38.485 154.570 ;
        RECT 40.050 154.305 42.745 154.570 ;
        RECT 5.240 153.690 42.745 154.305 ;
        RECT 5.240 153.490 5.590 153.690 ;
        RECT 9.865 153.490 10.265 153.540 ;
        RECT 8.340 153.290 10.265 153.490 ;
        RECT 8.340 142.365 8.540 153.290 ;
        RECT 9.865 153.240 10.265 153.290 ;
        RECT 18.565 152.740 18.865 153.140 ;
        RECT 29.340 152.740 31.040 153.690 ;
        RECT 36.590 152.890 36.890 153.290 ;
        RECT 18.565 143.565 18.765 152.740 ;
        RECT 23.640 152.290 23.940 152.690 ;
        RECT 18.565 143.140 18.815 143.565 ;
        RECT 18.615 142.365 18.815 143.140 ;
        RECT 23.690 142.365 23.890 152.290 ;
        RECT 26.240 151.840 26.540 152.240 ;
        RECT 26.290 142.365 26.490 151.840 ;
        RECT 27.490 151.390 27.790 151.790 ;
        RECT 27.540 142.365 27.740 151.390 ;
        RECT 28.690 150.940 28.990 151.340 ;
        RECT 28.740 142.365 28.940 150.940 ;
        RECT 29.940 150.490 30.240 150.890 ;
        RECT 29.990 142.365 30.190 150.490 ;
        RECT 31.140 150.040 31.440 150.440 ;
        RECT 31.190 142.365 31.390 150.040 ;
        RECT 32.340 149.590 32.640 149.990 ;
        RECT 32.390 142.365 32.590 149.590 ;
        RECT 33.590 149.140 33.890 149.540 ;
        RECT 33.640 142.365 33.840 149.140 ;
        RECT 34.740 148.690 35.040 149.090 ;
        RECT 34.790 142.365 34.990 148.690 ;
        RECT 36.640 146.840 36.840 152.890 ;
        RECT 44.135 150.380 44.635 154.980 ;
        RECT 55.485 150.430 55.985 154.980 ;
        RECT 61.435 150.430 61.935 154.980 ;
        RECT 70.235 150.430 70.735 154.980 ;
        RECT 43.885 149.980 44.685 150.380 ;
        RECT 55.285 150.130 56.035 150.430 ;
        RECT 55.285 149.980 55.585 150.130 ;
        RECT 55.735 149.980 56.035 150.130 ;
        RECT 61.185 150.180 61.935 150.430 ;
        RECT 61.185 149.980 61.485 150.180 ;
        RECT 61.635 149.980 61.935 150.180 ;
        RECT 70.135 150.180 70.885 150.430 ;
        RECT 70.135 149.980 70.435 150.180 ;
        RECT 70.585 149.980 70.885 150.180 ;
        RECT 47.340 148.690 47.640 149.090 ;
        RECT 37.490 148.240 37.790 148.640 ;
        RECT 36.590 146.440 36.890 146.840 ;
        RECT 8.240 141.965 8.640 142.365 ;
        RECT 18.540 141.965 18.840 142.365 ;
        RECT 23.640 141.965 23.940 142.365 ;
        RECT 26.240 141.965 26.540 142.365 ;
        RECT 27.490 141.965 27.790 142.365 ;
        RECT 28.690 141.965 28.990 142.365 ;
        RECT 29.940 141.965 30.240 142.365 ;
        RECT 31.140 141.965 31.440 142.365 ;
        RECT 32.340 141.965 32.640 142.365 ;
        RECT 33.590 141.965 33.890 142.365 ;
        RECT 34.740 141.965 35.040 142.365 ;
        RECT 37.540 142.265 37.740 148.240 ;
        RECT 41.340 147.790 41.640 148.190 ;
        RECT 41.390 142.265 41.590 147.790 ;
        RECT 43.290 147.340 43.590 147.740 ;
        RECT 43.340 142.265 43.540 147.340 ;
        RECT 44.140 146.890 44.440 147.290 ;
        RECT 44.190 142.265 44.390 146.890 ;
        RECT 45.240 146.440 45.540 146.840 ;
        RECT 45.290 142.265 45.490 146.440 ;
        RECT 47.390 142.265 47.590 148.690 ;
        RECT 51.190 148.240 51.490 148.640 ;
        RECT 51.240 142.265 51.440 148.240 ;
        RECT 55.040 147.790 55.340 148.190 ;
        RECT 55.090 142.265 55.290 147.790 ;
        RECT 56.940 147.340 57.240 147.740 ;
        RECT 56.990 142.265 57.190 147.340 ;
        RECT 57.890 146.890 58.190 147.290 ;
        RECT 57.940 142.265 58.140 146.890 ;
        RECT 65.340 146.440 65.640 146.840 ;
        RECT 58.940 145.990 59.240 146.390 ;
        RECT 58.990 142.265 59.190 145.990 ;
        RECT 59.890 145.540 60.190 145.940 ;
        RECT 59.940 142.265 60.140 145.540 ;
        RECT 60.490 145.090 60.790 145.490 ;
        RECT 60.540 142.265 60.740 145.090 ;
        RECT 61.540 144.640 61.840 145.040 ;
        RECT 61.590 142.265 61.790 144.640 ;
        RECT 62.590 144.190 62.890 144.590 ;
        RECT 62.640 142.265 62.840 144.190 ;
        RECT 63.640 143.740 63.940 144.140 ;
        RECT 63.690 142.265 63.890 143.740 ;
        RECT 64.690 143.290 64.990 143.690 ;
        RECT 64.740 142.265 64.940 143.290 ;
        RECT 37.490 141.865 37.790 142.265 ;
        RECT 41.340 141.865 41.640 142.265 ;
        RECT 43.290 141.865 43.590 142.265 ;
        RECT 44.140 141.865 44.440 142.265 ;
        RECT 45.240 141.865 45.540 142.265 ;
        RECT 47.340 141.865 47.640 142.265 ;
        RECT 51.190 141.865 51.490 142.265 ;
        RECT 55.040 141.865 55.340 142.265 ;
        RECT 56.940 141.865 57.240 142.265 ;
        RECT 57.890 141.865 58.190 142.265 ;
        RECT 58.940 141.865 59.240 142.265 ;
        RECT 59.890 141.865 60.190 142.265 ;
        RECT 60.490 141.865 60.790 142.265 ;
        RECT 61.540 141.865 61.840 142.265 ;
        RECT 62.590 141.865 62.890 142.265 ;
        RECT 63.640 141.865 63.940 142.265 ;
        RECT 64.690 141.865 64.990 142.265 ;
        RECT 5.890 141.565 6.190 141.640 ;
        RECT 46.640 141.565 46.940 141.665 ;
        RECT 47.590 141.565 47.890 141.665 ;
        RECT 48.540 141.565 48.840 141.665 ;
        RECT 49.490 141.565 49.790 141.665 ;
        RECT 50.490 141.565 50.790 141.665 ;
        RECT 51.440 141.565 51.740 141.665 ;
        RECT 52.390 141.565 52.690 141.665 ;
        RECT 53.340 141.565 53.640 141.665 ;
        RECT 54.340 141.565 54.640 141.665 ;
        RECT 55.290 141.565 55.590 141.665 ;
        RECT 56.240 141.565 56.540 141.665 ;
        RECT 57.190 141.565 57.490 141.665 ;
        RECT 5.890 141.365 57.490 141.565 ;
        RECT 5.890 141.240 6.190 141.365 ;
        RECT 46.640 141.265 46.940 141.365 ;
        RECT 47.590 141.265 47.890 141.365 ;
        RECT 48.540 141.265 48.840 141.365 ;
        RECT 49.490 141.265 49.790 141.365 ;
        RECT 50.490 141.265 50.790 141.365 ;
        RECT 51.440 141.265 51.740 141.365 ;
        RECT 52.390 141.265 52.690 141.365 ;
        RECT 53.340 141.265 53.640 141.365 ;
        RECT 54.340 141.265 54.640 141.365 ;
        RECT 55.290 141.265 55.590 141.365 ;
        RECT 56.240 141.215 56.540 141.365 ;
        RECT 57.190 141.265 57.490 141.365 ;
        RECT 58.240 141.065 58.540 141.165 ;
        RECT 59.190 141.065 59.490 141.165 ;
        RECT 60.240 141.065 60.540 141.165 ;
        RECT 61.290 141.065 61.590 141.165 ;
        RECT 62.340 141.065 62.640 141.165 ;
        RECT 63.390 141.065 63.690 141.165 ;
        RECT 64.440 141.065 64.740 141.165 ;
        RECT 5.240 140.065 5.540 140.140 ;
        RECT 7.340 140.065 7.640 140.915 ;
        RECT 57.190 140.865 64.740 141.065 ;
        RECT 57.190 140.815 58.540 140.865 ;
        RECT 57.190 140.665 57.490 140.815 ;
        RECT 58.290 140.765 58.540 140.815 ;
        RECT 59.190 140.765 59.490 140.865 ;
        RECT 60.240 140.765 60.540 140.865 ;
        RECT 61.290 140.765 61.590 140.865 ;
        RECT 62.340 140.765 62.640 140.865 ;
        RECT 63.390 140.765 63.690 140.865 ;
        RECT 64.440 140.765 64.740 140.865 ;
        RECT 47.140 140.565 47.440 140.665 ;
        RECT 48.090 140.565 48.390 140.665 ;
        RECT 48.590 140.565 48.890 140.665 ;
        RECT 49.040 140.565 49.340 140.665 ;
        RECT 49.990 140.565 50.290 140.665 ;
        RECT 47.140 140.365 50.290 140.565 ;
        RECT 47.140 140.265 47.440 140.365 ;
        RECT 48.090 140.265 48.390 140.365 ;
        RECT 48.590 140.265 48.890 140.365 ;
        RECT 49.040 140.265 49.340 140.365 ;
        RECT 49.990 140.265 50.290 140.365 ;
        RECT 5.240 139.865 7.640 140.065 ;
        RECT 5.240 139.740 5.540 139.865 ;
        RECT 7.340 139.015 7.640 139.865 ;
        RECT 4.590 138.515 4.890 138.590 ;
        RECT 7.940 138.515 8.240 138.615 ;
        RECT 9.240 138.515 9.540 138.615 ;
        RECT 10.540 138.515 10.840 138.615 ;
        RECT 11.790 138.515 12.090 138.615 ;
        RECT 13.090 138.515 13.390 138.615 ;
        RECT 14.340 138.515 14.640 138.615 ;
        RECT 15.640 138.515 15.940 138.615 ;
        RECT 16.940 138.515 17.240 138.615 ;
        RECT 18.190 138.515 18.490 138.615 ;
        RECT 19.490 138.515 19.790 138.615 ;
        RECT 20.740 138.515 21.040 138.615 ;
        RECT 22.040 138.515 22.340 138.615 ;
        RECT 23.340 138.515 23.640 138.615 ;
        RECT 24.590 138.515 24.890 138.615 ;
        RECT 25.890 138.515 26.190 138.615 ;
        RECT 27.190 138.515 27.490 138.615 ;
        RECT 28.390 138.515 28.690 138.615 ;
        RECT 29.590 138.515 29.890 138.615 ;
        RECT 30.790 138.515 31.090 138.615 ;
        RECT 32.040 138.515 32.340 138.615 ;
        RECT 33.240 138.515 33.540 138.615 ;
        RECT 34.440 138.515 34.740 138.615 ;
        RECT 4.590 138.315 34.740 138.515 ;
        RECT 4.590 138.190 4.890 138.315 ;
        RECT 7.940 138.215 8.240 138.315 ;
        RECT 9.240 138.215 9.540 138.315 ;
        RECT 10.540 138.215 10.840 138.315 ;
        RECT 11.790 138.215 12.090 138.315 ;
        RECT 13.090 138.215 13.390 138.315 ;
        RECT 14.340 138.215 14.640 138.315 ;
        RECT 15.640 138.215 15.940 138.315 ;
        RECT 16.940 138.215 17.240 138.315 ;
        RECT 18.190 138.215 18.490 138.315 ;
        RECT 19.490 138.215 19.790 138.315 ;
        RECT 20.740 138.215 21.040 138.315 ;
        RECT 22.040 138.215 22.340 138.315 ;
        RECT 23.340 138.215 23.640 138.315 ;
        RECT 24.590 138.215 24.890 138.315 ;
        RECT 25.890 138.215 26.190 138.315 ;
        RECT 27.190 138.215 27.490 138.315 ;
        RECT 28.390 138.215 28.690 138.315 ;
        RECT 29.590 138.215 29.890 138.315 ;
        RECT 30.790 138.215 31.090 138.315 ;
        RECT 32.040 138.215 32.340 138.315 ;
        RECT 33.240 138.215 33.540 138.315 ;
        RECT 34.440 138.215 34.740 138.315 ;
        RECT 35.290 138.240 36.990 140.040 ;
        RECT 58.740 139.915 59.040 140.315 ;
        RECT 59.690 139.915 59.990 140.315 ;
        RECT 60.740 139.915 61.040 140.315 ;
        RECT 61.790 139.915 62.090 140.315 ;
        RECT 62.840 139.915 63.140 140.315 ;
        RECT 63.890 139.965 64.190 140.365 ;
        RECT 64.940 139.965 65.240 140.365 ;
        RECT 45.240 139.515 45.540 139.615 ;
        RECT 64.190 139.515 64.490 139.615 ;
        RECT 45.240 139.315 64.490 139.515 ;
        RECT 45.240 139.215 45.540 139.315 ;
        RECT 64.190 139.215 64.490 139.315 ;
        RECT 58.990 138.765 59.290 139.165 ;
        RECT 43.490 138.365 43.790 138.465 ;
        RECT 57.190 138.365 57.490 138.465 ;
        RECT 43.490 138.165 57.490 138.365 ;
        RECT 43.490 138.065 43.790 138.165 ;
        RECT 57.190 138.065 57.490 138.165 ;
        RECT 3.940 136.465 4.240 136.540 ;
        RECT 36.790 136.465 37.090 136.565 ;
        RECT 37.740 136.465 38.040 136.565 ;
        RECT 38.690 136.465 38.990 136.565 ;
        RECT 39.690 136.465 39.990 136.565 ;
        RECT 40.640 136.465 40.940 136.565 ;
        RECT 41.590 136.465 41.890 136.565 ;
        RECT 42.540 136.465 42.840 136.565 ;
        RECT 43.490 136.465 43.790 136.565 ;
        RECT 3.940 136.265 43.790 136.465 ;
        RECT 59.040 136.265 59.240 138.765 ;
        RECT 59.940 138.415 60.240 138.815 ;
        RECT 59.990 136.265 60.190 138.415 ;
        RECT 60.490 138.015 60.790 138.415 ;
        RECT 60.540 136.265 60.740 138.015 ;
        RECT 61.540 137.615 61.840 138.015 ;
        RECT 61.590 136.265 61.790 137.615 ;
        RECT 62.590 137.215 62.890 137.615 ;
        RECT 62.640 136.265 62.840 137.215 ;
        RECT 63.640 136.815 63.940 137.215 ;
        RECT 65.390 136.815 65.590 146.440 ;
        RECT 66.140 145.990 66.440 146.390 ;
        RECT 65.740 144.640 66.040 145.040 ;
        RECT 63.690 136.265 63.890 136.815 ;
        RECT 64.690 136.415 64.990 136.815 ;
        RECT 65.340 136.415 65.640 136.815 ;
        RECT 64.740 136.265 64.940 136.415 ;
        RECT 65.790 136.265 65.990 144.640 ;
        RECT 66.190 137.215 66.390 145.990 ;
        RECT 66.940 145.540 67.240 145.940 ;
        RECT 66.540 144.190 66.840 144.590 ;
        RECT 66.590 138.415 66.790 144.190 ;
        RECT 66.540 138.015 66.840 138.415 ;
        RECT 66.990 137.615 67.190 145.540 ;
        RECT 67.740 145.090 68.040 145.490 ;
        RECT 67.340 143.740 67.640 144.140 ;
        RECT 67.390 138.815 67.590 143.740 ;
        RECT 67.340 138.415 67.640 138.815 ;
        RECT 67.790 138.015 67.990 145.090 ;
        RECT 77.615 143.690 77.765 161.340 ;
        RECT 78.065 144.140 78.215 161.640 ;
        RECT 78.515 144.590 78.665 161.940 ;
        RECT 78.965 145.040 79.115 162.240 ;
        RECT 79.415 145.490 79.565 162.540 ;
        RECT 79.865 145.940 80.015 162.840 ;
        RECT 80.315 163.140 80.615 163.540 ;
        RECT 80.315 146.390 80.465 163.140 ;
        RECT 80.765 162.840 81.065 163.240 ;
        RECT 80.765 146.840 80.915 162.840 ;
        RECT 81.215 162.540 81.515 162.940 ;
        RECT 81.215 147.290 81.365 162.540 ;
        RECT 81.665 162.240 81.965 162.640 ;
        RECT 81.665 147.740 81.815 162.240 ;
        RECT 82.115 161.940 82.415 162.340 ;
        RECT 82.115 148.190 82.265 161.940 ;
        RECT 82.565 161.640 82.865 162.040 ;
        RECT 82.565 148.640 82.715 161.640 ;
        RECT 83.015 161.340 83.315 161.740 ;
        RECT 83.015 149.090 83.165 161.340 ;
        RECT 105.340 161.290 105.490 163.640 ;
        RECT 125.195 162.065 125.495 169.365 ;
        RECT 138.745 164.015 138.945 169.365 ;
        RECT 142.385 169.265 142.685 169.365 ;
        RECT 142.925 169.515 143.225 169.665 ;
        RECT 145.295 169.515 145.595 169.665 ;
        RECT 142.925 169.365 145.595 169.515 ;
        RECT 142.925 169.265 143.225 169.365 ;
        RECT 145.295 169.265 145.595 169.365 ;
        RECT 142.645 168.965 142.995 169.115 ;
        RECT 145.845 168.965 146.145 169.065 ;
        RECT 142.645 168.765 146.145 168.965 ;
        RECT 139.445 168.365 139.745 168.765 ;
        RECT 142.645 168.665 142.995 168.765 ;
        RECT 145.845 168.665 146.145 168.765 ;
        RECT 139.495 166.015 139.695 168.365 ;
        RECT 143.595 168.015 143.895 168.165 ;
        RECT 146.195 168.015 146.495 168.165 ;
        RECT 143.595 167.865 146.495 168.015 ;
        RECT 143.595 167.765 143.895 167.865 ;
        RECT 146.195 167.765 146.495 167.865 ;
        RECT 142.045 167.615 142.345 167.715 ;
        RECT 144.445 167.615 144.745 167.715 ;
        RECT 148.895 167.615 149.195 167.715 ;
        RECT 142.045 167.415 149.195 167.615 ;
        RECT 142.045 167.315 142.345 167.415 ;
        RECT 144.445 167.315 144.745 167.415 ;
        RECT 148.895 167.315 149.195 167.415 ;
        RECT 143.695 167.115 143.995 167.215 ;
        RECT 146.695 167.115 146.995 167.265 ;
        RECT 143.695 166.965 146.995 167.115 ;
        RECT 143.695 166.815 143.995 166.965 ;
        RECT 146.695 166.865 146.995 166.965 ;
        RECT 142.745 166.665 143.045 166.715 ;
        RECT 145.845 166.665 146.145 166.815 ;
        RECT 148.345 166.665 148.645 166.765 ;
        RECT 142.745 166.515 148.645 166.665 ;
        RECT 142.745 166.315 143.045 166.515 ;
        RECT 145.845 166.415 146.145 166.515 ;
        RECT 148.345 166.365 148.645 166.515 ;
        RECT 142.440 166.015 142.740 166.135 ;
        RECT 139.495 165.815 142.740 166.015 ;
        RECT 142.440 165.735 142.740 165.815 ;
        RECT 142.980 166.015 143.280 166.135 ;
        RECT 144.995 166.015 145.295 166.115 ;
        RECT 142.980 165.865 145.295 166.015 ;
        RECT 142.980 165.735 143.280 165.865 ;
        RECT 144.995 165.715 145.295 165.865 ;
        RECT 143.195 165.015 143.495 165.165 ;
        RECT 147.145 165.015 147.445 165.115 ;
        RECT 143.195 164.865 147.445 165.015 ;
        RECT 143.195 164.765 143.495 164.865 ;
        RECT 147.145 164.715 147.445 164.865 ;
        RECT 142.440 164.015 142.740 164.135 ;
        RECT 138.745 163.815 142.740 164.015 ;
        RECT 142.440 163.735 142.740 163.815 ;
        RECT 142.980 164.065 143.280 164.135 ;
        RECT 145.395 164.065 145.695 164.165 ;
        RECT 142.980 163.865 145.695 164.065 ;
        RECT 142.980 163.735 143.280 163.865 ;
        RECT 145.395 163.765 145.695 163.865 ;
        RECT 142.695 163.365 142.995 163.565 ;
        RECT 145.845 163.365 146.145 163.615 ;
        RECT 142.695 163.215 146.145 163.365 ;
        RECT 142.695 163.165 142.995 163.215 ;
        RECT 143.645 162.815 143.945 162.915 ;
        RECT 146.145 162.815 146.445 162.915 ;
        RECT 143.645 162.665 146.445 162.815 ;
        RECT 143.645 162.515 143.945 162.665 ;
        RECT 146.145 162.515 146.445 162.665 ;
        RECT 105.240 160.890 105.540 161.290 ;
        RECT 128.890 160.245 130.590 160.290 ;
        RECT 123.565 159.780 140.910 160.245 ;
        RECT 128.890 159.740 130.590 159.780 ;
        RECT 90.195 159.240 91.070 159.500 ;
        RECT 99.055 159.240 99.930 159.500 ;
        RECT 104.955 159.240 105.830 159.500 ;
        RECT 116.335 159.250 117.210 159.510 ;
        RECT 118.845 159.505 119.720 159.565 ;
        RECT 133.195 159.505 134.070 159.610 ;
        RECT 118.845 159.350 134.070 159.505 ;
        RECT 118.845 159.345 133.195 159.350 ;
        RECT 118.845 159.305 119.720 159.345 ;
        RECT 90.380 155.240 90.880 159.240 ;
        RECT 99.180 155.240 99.680 159.240 ;
        RECT 105.130 155.240 105.630 159.240 ;
        RECT 116.480 156.630 116.980 159.250 ;
        RECT 119.960 157.360 120.120 159.345 ;
        RECT 138.615 158.895 139.615 159.780 ;
        RECT 129.180 158.810 137.920 158.870 ;
        RECT 120.515 158.420 120.775 158.700 ;
        RECT 121.475 158.420 121.735 158.700 ;
        RECT 122.435 158.420 122.695 158.700 ;
        RECT 120.515 158.160 122.695 158.420 ;
        RECT 120.515 157.825 120.775 158.160 ;
        RECT 121.475 157.825 121.735 158.160 ;
        RECT 122.435 157.825 122.695 158.160 ;
        RECT 129.175 158.610 137.920 158.810 ;
        RECT 140.175 158.790 141.175 159.235 ;
        RECT 150.525 158.840 150.825 158.890 ;
        RECT 150.450 158.790 150.825 158.840 ;
        RECT 129.175 157.935 129.435 158.610 ;
        RECT 140.175 158.590 150.825 158.790 ;
        RECT 133.150 158.275 134.150 158.330 ;
        RECT 121.035 157.390 121.295 157.670 ;
        RECT 121.995 157.390 122.255 157.670 ;
        RECT 123.830 157.390 124.830 157.930 ;
        RECT 133.005 157.890 134.255 158.275 ;
        RECT 140.175 158.235 141.175 158.590 ;
        RECT 150.450 158.540 150.825 158.590 ;
        RECT 150.525 158.490 150.825 158.540 ;
        RECT 157.525 157.890 157.825 157.990 ;
        RECT 126.645 157.390 126.905 157.830 ;
        RECT 127.985 157.390 128.245 157.820 ;
        RECT 133.005 157.690 157.825 157.890 ;
        RECT 133.005 157.400 134.255 157.690 ;
        RECT 157.525 157.590 157.825 157.690 ;
        RECT 121.035 157.360 128.245 157.390 ;
        RECT 119.960 157.200 128.245 157.360 ;
        RECT 133.150 157.330 134.150 157.400 ;
        RECT 121.035 157.130 128.245 157.200 ;
        RECT 121.035 156.795 121.295 157.130 ;
        RECT 121.995 156.795 122.255 157.130 ;
        RECT 123.830 156.930 124.830 157.130 ;
        RECT 126.645 156.955 126.905 157.130 ;
        RECT 127.985 156.945 128.245 157.130 ;
        RECT 133.525 156.630 133.785 157.010 ;
        RECT 135.575 156.630 135.835 157.060 ;
        RECT 137.525 156.990 140.445 157.460 ;
        RECT 116.480 156.380 135.835 156.630 ;
        RECT 116.480 155.240 116.980 156.380 ;
        RECT 90.205 154.980 91.080 155.240 ;
        RECT 99.105 154.980 99.980 155.240 ;
        RECT 105.005 154.980 105.880 155.240 ;
        RECT 116.355 154.980 117.230 155.240 ;
        RECT 119.475 155.085 119.735 155.960 ;
        RECT 125.455 155.850 125.715 156.190 ;
        RECT 131.375 155.850 131.635 156.190 ;
        RECT 133.525 156.135 133.785 156.380 ;
        RECT 135.575 156.185 135.835 156.380 ;
        RECT 125.455 155.610 131.635 155.850 ;
        RECT 125.455 155.315 125.715 155.610 ;
        RECT 131.375 155.315 131.635 155.610 ;
        RECT 90.380 150.430 90.880 154.980 ;
        RECT 99.180 150.430 99.680 154.980 ;
        RECT 105.130 150.430 105.630 154.980 ;
        RECT 90.230 150.180 90.980 150.430 ;
        RECT 90.230 149.980 90.530 150.180 ;
        RECT 90.680 149.980 90.980 150.180 ;
        RECT 99.180 150.180 99.930 150.430 ;
        RECT 99.180 149.980 99.480 150.180 ;
        RECT 99.630 149.980 99.930 150.180 ;
        RECT 105.080 150.130 105.830 150.430 ;
        RECT 116.480 150.380 116.980 154.980 ;
        RECT 119.530 154.570 119.680 155.085 ;
        RECT 124.115 154.980 131.170 155.165 ;
        RECT 137.340 155.155 137.600 156.030 ;
        RECT 138.705 155.240 139.705 156.240 ;
        RECT 137.380 154.980 137.530 155.155 ;
        RECT 121.250 154.965 137.530 154.980 ;
        RECT 121.250 154.780 124.360 154.965 ;
        RECT 130.930 154.780 137.530 154.965 ;
        RECT 121.250 154.665 122.255 154.780 ;
        RECT 130.930 154.710 131.995 154.780 ;
        RECT 135.305 154.710 136.180 154.780 ;
        RECT 125.160 154.570 126.035 154.675 ;
        RECT 128.485 154.570 129.360 154.675 ;
        RECT 138.450 154.570 139.450 154.695 ;
        RECT 139.990 154.570 140.445 156.990 ;
        RECT 155.525 154.570 155.875 154.790 ;
        RECT 118.370 154.305 121.065 154.570 ;
        RECT 122.630 154.305 155.875 154.570 ;
        RECT 118.370 153.690 155.875 154.305 ;
        RECT 124.225 152.890 124.525 153.290 ;
        RECT 105.080 149.980 105.380 150.130 ;
        RECT 105.530 149.980 105.830 150.130 ;
        RECT 116.430 149.980 117.230 150.380 ;
        RECT 82.940 148.690 83.240 149.090 ;
        RECT 113.475 148.690 113.775 149.090 ;
        RECT 82.490 148.240 82.790 148.640 ;
        RECT 109.625 148.240 109.925 148.640 ;
        RECT 82.040 147.790 82.340 148.190 ;
        RECT 105.775 147.790 106.075 148.190 ;
        RECT 81.590 147.340 81.890 147.740 ;
        RECT 103.875 147.340 104.175 147.740 ;
        RECT 81.140 146.890 81.440 147.290 ;
        RECT 102.925 146.890 103.225 147.290 ;
        RECT 80.690 146.440 80.990 146.840 ;
        RECT 95.475 146.440 95.775 146.840 ;
        RECT 80.240 145.990 80.540 146.390 ;
        RECT 94.675 145.990 94.975 146.390 ;
        RECT 79.790 145.540 80.090 145.940 ;
        RECT 93.875 145.540 94.175 145.940 ;
        RECT 79.340 145.090 79.640 145.490 ;
        RECT 93.075 145.090 93.375 145.490 ;
        RECT 78.890 144.640 79.190 145.040 ;
        RECT 78.440 144.190 78.740 144.590 ;
        RECT 77.990 143.740 78.290 144.140 ;
        RECT 68.140 143.290 68.440 143.690 ;
        RECT 77.540 143.290 77.840 143.690 ;
        RECT 92.675 143.290 92.975 143.690 ;
        RECT 68.190 139.215 68.390 143.290 ;
        RECT 72.690 141.215 72.990 141.615 ;
        RECT 72.740 139.565 72.890 141.215 ;
        RECT 74.490 141.015 74.790 141.415 ;
        RECT 86.325 141.015 86.625 141.415 ;
        RECT 88.125 141.215 88.425 141.615 ;
        RECT 68.140 138.815 68.440 139.215 ;
        RECT 72.690 139.165 72.990 139.565 ;
        RECT 67.740 137.615 68.040 138.015 ;
        RECT 66.940 137.215 67.240 137.615 ;
        RECT 72.740 137.415 72.890 139.165 ;
        RECT 74.090 139.015 74.390 139.415 ;
        RECT 66.140 136.815 66.440 137.215 ;
        RECT 72.690 137.015 72.990 137.415 ;
        RECT 3.940 136.140 4.240 136.265 ;
        RECT 36.790 136.165 37.090 136.265 ;
        RECT 37.740 136.165 38.040 136.265 ;
        RECT 38.690 136.165 38.990 136.265 ;
        RECT 39.690 136.165 39.990 136.265 ;
        RECT 40.640 136.165 40.940 136.265 ;
        RECT 41.590 136.165 41.890 136.265 ;
        RECT 42.540 136.165 42.840 136.265 ;
        RECT 43.490 136.165 43.790 136.265 ;
        RECT 3.290 135.815 3.590 135.890 ;
        RECT 44.540 135.815 44.840 135.915 ;
        RECT 45.490 135.815 45.790 135.915 ;
        RECT 58.990 135.865 59.290 136.265 ;
        RECT 59.940 135.865 60.240 136.265 ;
        RECT 60.490 135.865 60.790 136.265 ;
        RECT 61.540 135.865 61.840 136.265 ;
        RECT 62.590 135.865 62.890 136.265 ;
        RECT 63.640 135.865 63.940 136.265 ;
        RECT 64.690 135.865 64.990 136.265 ;
        RECT 65.740 135.865 66.040 136.265 ;
        RECT 3.290 135.615 45.790 135.815 ;
        RECT 3.290 135.490 3.590 135.615 ;
        RECT 44.540 135.515 44.840 135.615 ;
        RECT 45.465 135.515 45.790 135.615 ;
        RECT 56.240 135.665 56.540 135.715 ;
        RECT 58.240 135.665 58.540 135.715 ;
        RECT 59.190 135.665 59.490 135.715 ;
        RECT 60.240 135.665 60.540 135.715 ;
        RECT 61.290 135.665 61.590 135.715 ;
        RECT 62.340 135.665 62.640 135.715 ;
        RECT 63.390 135.665 63.690 135.715 ;
        RECT 64.440 135.665 64.740 135.715 ;
        RECT 65.490 135.665 65.790 135.715 ;
        RECT 45.465 134.965 45.715 135.515 ;
        RECT 56.240 135.365 65.790 135.665 ;
        RECT 56.240 135.315 56.540 135.365 ;
        RECT 58.240 135.315 58.540 135.365 ;
        RECT 59.190 135.315 59.490 135.365 ;
        RECT 60.240 135.315 60.540 135.365 ;
        RECT 61.290 135.315 61.590 135.365 ;
        RECT 62.340 135.315 62.640 135.365 ;
        RECT 63.390 135.315 63.690 135.365 ;
        RECT 64.440 135.315 64.740 135.365 ;
        RECT 65.490 135.315 65.790 135.365 ;
        RECT 66.540 135.615 66.840 135.715 ;
        RECT 67.490 135.615 67.790 135.715 ;
        RECT 69.040 135.615 69.340 135.715 ;
        RECT 70.090 135.615 70.390 135.715 ;
        RECT 71.140 135.615 71.440 135.715 ;
        RECT 72.190 135.615 72.490 135.715 ;
        RECT 72.740 135.615 72.890 137.015 ;
        RECT 73.690 136.765 73.990 137.165 ;
        RECT 73.240 135.615 73.540 135.715 ;
        RECT 66.540 135.415 73.540 135.615 ;
        RECT 66.540 135.315 66.840 135.415 ;
        RECT 67.490 135.315 67.790 135.415 ;
        RECT 69.040 135.315 69.340 135.415 ;
        RECT 70.090 135.315 70.390 135.415 ;
        RECT 71.140 135.315 71.440 135.415 ;
        RECT 72.190 135.315 72.490 135.415 ;
        RECT 73.240 135.315 73.540 135.415 ;
        RECT 66.640 134.965 66.790 135.315 ;
        RECT 45.465 134.715 66.790 134.965 ;
        RECT 68.540 134.765 68.840 135.165 ;
        RECT 69.590 134.765 69.890 135.165 ;
        RECT 70.640 134.765 70.940 135.165 ;
        RECT 71.690 134.765 71.990 135.165 ;
        RECT 72.740 134.765 73.040 135.165 ;
        RECT 37.290 134.265 37.590 134.365 ;
        RECT 38.240 134.265 38.540 134.365 ;
        RECT 39.190 134.265 39.490 134.365 ;
        RECT 40.140 134.265 40.440 134.365 ;
        RECT 8.590 134.165 8.890 134.265 ;
        RECT 9.890 134.165 10.190 134.265 ;
        RECT 11.190 134.165 11.490 134.265 ;
        RECT 12.440 134.165 12.740 134.265 ;
        RECT 13.740 134.165 14.040 134.265 ;
        RECT 14.990 134.165 15.290 134.265 ;
        RECT 16.290 134.165 16.590 134.265 ;
        RECT 17.590 134.165 17.890 134.265 ;
        RECT 8.590 133.965 17.890 134.165 ;
        RECT 8.590 133.865 8.890 133.965 ;
        RECT 9.890 133.865 10.190 133.965 ;
        RECT 11.190 133.865 11.490 133.965 ;
        RECT 12.440 133.865 12.740 133.965 ;
        RECT 13.740 133.865 14.040 133.965 ;
        RECT 14.990 133.865 15.290 133.965 ;
        RECT 16.290 133.865 16.590 133.965 ;
        RECT 17.590 133.865 17.890 133.965 ;
        RECT 18.840 134.165 19.140 134.265 ;
        RECT 20.140 134.165 20.440 134.265 ;
        RECT 21.390 134.165 21.690 134.265 ;
        RECT 22.690 134.165 22.990 134.265 ;
        RECT 18.840 133.965 22.990 134.165 ;
        RECT 18.840 133.865 19.140 133.965 ;
        RECT 20.140 133.865 20.440 133.965 ;
        RECT 21.390 133.865 21.690 133.965 ;
        RECT 22.690 133.865 22.990 133.965 ;
        RECT 23.940 134.165 24.240 134.265 ;
        RECT 25.240 134.165 25.540 134.265 ;
        RECT 23.940 133.965 25.540 134.165 ;
        RECT 23.940 133.865 24.240 133.965 ;
        RECT 25.240 133.865 25.540 133.965 ;
        RECT 26.540 133.865 26.840 134.265 ;
        RECT 27.790 133.865 28.090 134.265 ;
        RECT 8.640 132.740 8.840 133.865 ;
        RECT 8.590 132.340 8.890 132.740 ;
        RECT 18.890 132.290 19.090 133.865 ;
        RECT 18.840 131.890 19.140 132.290 ;
        RECT 23.990 131.840 24.190 133.865 ;
        RECT 23.940 131.440 24.240 131.840 ;
        RECT 26.590 131.390 26.790 133.865 ;
        RECT 26.540 130.990 26.840 131.390 ;
        RECT 27.840 130.940 28.040 133.865 ;
        RECT 29.040 133.715 29.340 134.115 ;
        RECT 30.240 133.715 30.540 134.115 ;
        RECT 31.440 133.715 31.740 134.115 ;
        RECT 32.690 133.715 32.990 134.115 ;
        RECT 33.890 133.715 34.190 134.115 ;
        RECT 35.090 133.715 35.390 134.115 ;
        RECT 37.290 134.065 40.440 134.265 ;
        RECT 37.290 133.965 37.590 134.065 ;
        RECT 38.240 133.965 38.540 134.065 ;
        RECT 39.190 133.965 39.490 134.065 ;
        RECT 40.140 133.965 40.440 134.065 ;
        RECT 41.090 134.265 41.390 134.365 ;
        RECT 42.090 134.265 42.390 134.365 ;
        RECT 41.090 134.065 42.390 134.265 ;
        RECT 41.090 133.965 41.390 134.065 ;
        RECT 42.090 133.965 42.390 134.065 ;
        RECT 43.040 133.965 43.340 134.365 ;
        RECT 43.990 133.965 44.290 134.365 ;
        RECT 45.040 133.965 45.340 134.365 ;
        RECT 45.990 133.965 46.290 134.365 ;
        RECT 50.940 134.115 51.240 134.215 ;
        RECT 51.940 134.115 52.240 134.215 ;
        RECT 52.890 134.115 53.190 134.215 ;
        RECT 53.840 134.115 54.140 134.215 ;
        RECT 27.790 130.540 28.090 130.940 ;
        RECT 29.090 130.490 29.290 133.715 ;
        RECT 29.040 130.090 29.340 130.490 ;
        RECT 30.290 130.040 30.490 133.715 ;
        RECT 30.240 129.640 30.540 130.040 ;
        RECT 31.490 129.590 31.690 133.715 ;
        RECT 31.440 129.190 31.740 129.590 ;
        RECT 32.740 129.140 32.940 133.715 ;
        RECT 32.690 128.740 32.990 129.140 ;
        RECT 33.940 128.690 34.140 133.715 ;
        RECT 33.890 128.290 34.190 128.690 ;
        RECT 35.140 128.240 35.340 133.715 ;
        RECT 37.340 132.740 37.540 133.965 ;
        RECT 37.940 133.040 40.790 133.440 ;
        RECT 37.290 132.340 37.590 132.740 ;
        RECT 41.140 132.290 41.340 133.965 ;
        RECT 41.090 131.890 41.390 132.290 ;
        RECT 43.090 131.840 43.290 133.965 ;
        RECT 43.040 131.440 43.340 131.840 ;
        RECT 44.040 131.390 44.240 133.965 ;
        RECT 45.090 132.740 45.290 133.965 ;
        RECT 45.040 132.340 45.340 132.740 ;
        RECT 46.040 132.290 46.240 133.965 ;
        RECT 50.940 133.915 54.140 134.115 ;
        RECT 50.940 133.815 51.240 133.915 ;
        RECT 51.940 133.815 52.240 133.915 ;
        RECT 52.890 133.815 53.190 133.915 ;
        RECT 53.840 133.815 54.140 133.915 ;
        RECT 54.790 134.115 55.090 134.215 ;
        RECT 55.740 134.115 56.040 134.215 ;
        RECT 54.790 133.915 56.040 134.115 ;
        RECT 54.790 133.815 55.090 133.915 ;
        RECT 55.740 133.815 56.040 133.915 ;
        RECT 56.740 133.815 57.040 134.215 ;
        RECT 57.690 133.815 57.990 134.215 ;
        RECT 58.740 134.015 59.040 134.415 ;
        RECT 59.690 134.015 59.990 134.415 ;
        RECT 60.740 134.015 61.040 134.415 ;
        RECT 61.790 134.015 62.090 134.415 ;
        RECT 62.840 134.015 63.140 134.415 ;
        RECT 63.890 134.015 64.190 134.415 ;
        RECT 64.940 134.015 65.240 134.415 ;
        RECT 65.990 134.015 66.290 134.415 ;
        RECT 50.990 132.740 51.190 133.815 ;
        RECT 51.590 133.040 54.440 133.440 ;
        RECT 50.940 132.340 51.240 132.740 ;
        RECT 54.840 132.290 55.040 133.815 ;
        RECT 45.990 131.890 46.290 132.290 ;
        RECT 54.790 131.890 55.090 132.290 ;
        RECT 56.740 131.840 56.940 133.815 ;
        RECT 56.690 131.440 56.990 131.840 ;
        RECT 57.740 131.390 57.940 133.815 ;
        RECT 43.990 130.990 44.290 131.390 ;
        RECT 57.690 130.990 57.990 131.390 ;
        RECT 58.790 130.940 58.990 134.015 ;
        RECT 58.740 130.540 59.040 130.940 ;
        RECT 59.740 130.490 59.940 134.015 ;
        RECT 59.690 130.090 59.990 130.490 ;
        RECT 60.790 130.040 60.990 134.015 ;
        RECT 60.740 129.640 61.040 130.040 ;
        RECT 61.840 129.590 62.040 134.015 ;
        RECT 61.790 129.190 62.090 129.590 ;
        RECT 62.890 129.140 63.090 134.015 ;
        RECT 62.840 128.740 63.140 129.140 ;
        RECT 63.940 128.690 64.140 134.015 ;
        RECT 63.890 128.290 64.190 128.690 ;
        RECT 64.990 128.240 65.190 134.015 ;
        RECT 35.090 127.840 35.390 128.240 ;
        RECT 64.940 127.840 65.240 128.240 ;
        RECT 66.040 127.790 66.240 134.015 ;
        RECT 67.040 133.865 67.340 134.265 ;
        RECT 67.990 133.865 68.290 134.265 ;
        RECT 67.090 131.840 67.290 133.865 ;
        RECT 67.040 131.440 67.340 131.840 ;
        RECT 68.040 131.390 68.240 133.865 ;
        RECT 67.990 130.990 68.290 131.390 ;
        RECT 68.590 130.940 68.790 134.765 ;
        RECT 68.540 130.540 68.840 130.940 ;
        RECT 69.640 130.490 69.840 134.765 ;
        RECT 69.590 130.090 69.890 130.490 ;
        RECT 70.690 130.040 70.890 134.765 ;
        RECT 70.640 129.640 70.940 130.040 ;
        RECT 71.740 129.140 71.940 134.765 ;
        RECT 71.690 128.740 71.990 129.140 ;
        RECT 72.790 128.240 72.990 134.765 ;
        RECT 73.740 129.590 73.940 136.765 ;
        RECT 73.690 129.190 73.990 129.590 ;
        RECT 74.140 128.690 74.340 139.015 ;
        RECT 74.090 128.290 74.390 128.690 ;
        RECT 72.740 127.840 73.040 128.240 ;
        RECT 74.540 127.790 74.740 141.015 ;
        RECT 74.990 132.340 75.290 132.740 ;
        RECT 85.825 132.340 86.125 132.740 ;
        RECT 7.390 127.190 8.290 127.590 ;
        RECT 65.990 127.390 66.290 127.790 ;
        RECT 74.490 127.390 74.790 127.790 ;
        RECT 73.390 126.940 74.290 127.340 ;
        RECT 6.890 125.390 7.290 126.490 ;
        RECT 8.890 125.390 9.290 126.490 ;
        RECT 10.890 125.390 11.290 126.490 ;
        RECT 12.890 125.390 13.290 126.490 ;
        RECT 14.890 125.390 15.290 126.490 ;
        RECT 16.890 125.390 17.290 126.490 ;
        RECT 18.890 125.390 19.290 126.490 ;
        RECT 20.890 125.390 21.290 126.490 ;
        RECT 22.890 125.390 23.290 126.490 ;
        RECT 24.890 125.390 25.290 126.490 ;
        RECT 26.890 125.390 27.290 126.490 ;
        RECT 28.890 125.390 29.290 126.490 ;
        RECT 30.890 125.390 31.290 126.490 ;
        RECT 32.890 125.390 33.290 126.490 ;
        RECT 34.890 125.390 35.290 126.490 ;
        RECT 36.890 125.390 37.290 126.490 ;
        RECT 38.890 125.390 39.290 126.490 ;
        RECT 40.890 125.390 41.290 126.490 ;
        RECT 42.890 125.390 43.290 126.490 ;
        RECT 44.890 125.390 45.290 126.490 ;
        RECT 46.890 125.390 47.290 126.490 ;
        RECT 48.890 125.390 49.290 126.490 ;
        RECT 50.890 125.390 51.290 126.490 ;
        RECT 52.890 125.390 53.290 126.490 ;
        RECT 54.890 125.390 55.290 126.490 ;
        RECT 56.890 125.390 57.290 126.490 ;
        RECT 58.890 125.390 59.290 126.490 ;
        RECT 60.890 125.390 61.290 126.490 ;
        RECT 62.890 125.390 63.290 126.490 ;
        RECT 64.890 125.390 65.290 126.490 ;
        RECT 66.890 125.390 67.290 126.490 ;
        RECT 68.890 125.390 69.290 126.490 ;
        RECT 70.890 125.390 71.290 126.490 ;
        RECT 72.890 125.390 73.290 126.490 ;
        RECT 6.890 123.540 7.290 124.640 ;
        RECT 8.890 123.540 9.290 124.640 ;
        RECT 10.890 123.540 11.290 124.640 ;
        RECT 12.890 123.540 13.290 124.640 ;
        RECT 14.890 123.540 15.290 124.640 ;
        RECT 16.890 123.540 17.290 124.640 ;
        RECT 18.890 123.540 19.290 124.640 ;
        RECT 20.890 123.540 21.290 124.640 ;
        RECT 22.890 123.540 23.290 124.640 ;
        RECT 24.890 123.540 25.290 124.640 ;
        RECT 26.890 123.540 27.290 124.640 ;
        RECT 28.890 123.540 29.290 124.640 ;
        RECT 30.890 123.540 31.290 124.640 ;
        RECT 32.890 123.540 33.290 124.640 ;
        RECT 34.890 123.540 35.290 124.640 ;
        RECT 36.890 123.540 37.290 124.640 ;
        RECT 38.890 123.540 39.290 124.640 ;
        RECT 40.890 123.540 41.290 124.640 ;
        RECT 42.890 123.540 43.290 124.640 ;
        RECT 44.890 123.540 45.290 124.640 ;
        RECT 46.890 123.540 47.290 124.640 ;
        RECT 48.890 123.540 49.290 124.640 ;
        RECT 50.890 123.540 51.290 124.640 ;
        RECT 52.890 123.540 53.290 124.640 ;
        RECT 54.890 123.540 55.290 124.640 ;
        RECT 56.890 123.540 57.290 124.640 ;
        RECT 58.890 123.540 59.290 124.640 ;
        RECT 60.890 123.540 61.290 124.640 ;
        RECT 62.890 123.540 63.290 124.640 ;
        RECT 64.890 123.540 65.290 124.640 ;
        RECT 66.890 123.540 67.290 124.640 ;
        RECT 68.890 123.540 69.290 124.640 ;
        RECT 70.890 123.540 71.290 124.640 ;
        RECT 72.890 123.540 73.290 124.640 ;
        RECT 6.890 121.690 7.290 122.790 ;
        RECT 8.890 121.690 9.290 122.790 ;
        RECT 10.890 121.690 11.290 122.790 ;
        RECT 12.890 121.690 13.290 122.790 ;
        RECT 14.890 121.690 15.290 122.790 ;
        RECT 16.890 121.690 17.290 122.790 ;
        RECT 18.890 121.690 19.290 122.790 ;
        RECT 20.890 121.690 21.290 122.790 ;
        RECT 22.890 121.690 23.290 122.790 ;
        RECT 24.890 121.690 25.290 122.790 ;
        RECT 26.890 121.690 27.290 122.790 ;
        RECT 28.890 121.690 29.290 122.790 ;
        RECT 30.890 121.690 31.290 122.790 ;
        RECT 32.890 121.690 33.290 122.790 ;
        RECT 34.890 121.690 35.290 122.790 ;
        RECT 36.890 121.690 37.290 122.790 ;
        RECT 38.890 121.690 39.290 122.790 ;
        RECT 40.890 121.690 41.290 122.790 ;
        RECT 42.890 121.690 43.290 122.790 ;
        RECT 44.890 121.690 45.290 122.790 ;
        RECT 46.890 121.690 47.290 122.790 ;
        RECT 48.890 121.690 49.290 122.790 ;
        RECT 50.890 121.690 51.290 122.790 ;
        RECT 52.890 121.690 53.290 122.790 ;
        RECT 54.890 121.690 55.290 122.790 ;
        RECT 56.890 121.690 57.290 122.790 ;
        RECT 58.890 121.690 59.290 122.790 ;
        RECT 60.890 121.690 61.290 122.790 ;
        RECT 62.890 121.690 63.290 122.790 ;
        RECT 64.890 121.690 65.290 122.790 ;
        RECT 66.890 121.690 67.290 122.790 ;
        RECT 68.890 121.690 69.290 122.790 ;
        RECT 70.890 121.690 71.290 122.790 ;
        RECT 72.890 121.690 73.290 122.790 ;
        RECT 6.890 119.840 7.290 120.940 ;
        RECT 8.890 119.840 9.290 120.940 ;
        RECT 10.890 119.840 11.290 120.940 ;
        RECT 12.890 119.840 13.290 120.940 ;
        RECT 14.890 119.840 15.290 120.940 ;
        RECT 16.890 119.840 17.290 120.940 ;
        RECT 18.890 119.840 19.290 120.940 ;
        RECT 20.890 119.840 21.290 120.940 ;
        RECT 22.890 119.840 23.290 120.940 ;
        RECT 24.890 119.840 25.290 120.940 ;
        RECT 26.890 119.840 27.290 120.940 ;
        RECT 28.890 119.840 29.290 120.940 ;
        RECT 30.890 119.840 31.290 120.940 ;
        RECT 32.890 119.840 33.290 120.940 ;
        RECT 34.890 119.840 35.290 120.940 ;
        RECT 36.890 119.840 37.290 120.940 ;
        RECT 38.890 119.840 39.290 120.940 ;
        RECT 40.890 119.840 41.290 120.940 ;
        RECT 42.890 119.840 43.290 120.940 ;
        RECT 44.890 119.840 45.290 120.940 ;
        RECT 46.890 119.840 47.290 120.940 ;
        RECT 48.890 119.840 49.290 120.940 ;
        RECT 50.890 119.840 51.290 120.940 ;
        RECT 52.890 119.840 53.290 120.940 ;
        RECT 54.890 119.840 55.290 120.940 ;
        RECT 56.890 119.840 57.290 120.940 ;
        RECT 58.890 119.840 59.290 120.940 ;
        RECT 60.890 119.840 61.290 120.940 ;
        RECT 62.890 119.840 63.290 120.940 ;
        RECT 64.890 119.840 65.290 120.940 ;
        RECT 66.890 119.840 67.290 120.940 ;
        RECT 68.890 119.840 69.290 120.940 ;
        RECT 70.890 119.840 71.290 120.940 ;
        RECT 72.890 119.840 73.290 120.940 ;
        RECT 6.890 117.990 7.290 119.090 ;
        RECT 8.890 117.990 9.290 119.090 ;
        RECT 10.890 117.990 11.290 119.090 ;
        RECT 12.890 117.990 13.290 119.090 ;
        RECT 14.890 117.990 15.290 119.090 ;
        RECT 16.890 117.990 17.290 119.090 ;
        RECT 18.890 117.990 19.290 119.090 ;
        RECT 20.890 117.990 21.290 119.090 ;
        RECT 22.890 117.990 23.290 119.090 ;
        RECT 24.890 117.990 25.290 119.090 ;
        RECT 26.890 117.990 27.290 119.090 ;
        RECT 28.890 117.990 29.290 119.090 ;
        RECT 30.890 117.990 31.290 119.090 ;
        RECT 32.890 117.990 33.290 119.090 ;
        RECT 34.890 117.990 35.290 119.090 ;
        RECT 36.890 117.990 37.290 119.090 ;
        RECT 38.890 117.990 39.290 119.090 ;
        RECT 40.890 117.990 41.290 119.090 ;
        RECT 42.890 117.990 43.290 119.090 ;
        RECT 44.890 117.990 45.290 119.090 ;
        RECT 46.890 117.990 47.290 119.090 ;
        RECT 48.890 117.990 49.290 119.090 ;
        RECT 50.890 117.990 51.290 119.090 ;
        RECT 52.890 117.990 53.290 119.090 ;
        RECT 54.890 117.990 55.290 119.090 ;
        RECT 56.890 117.990 57.290 119.090 ;
        RECT 58.890 117.990 59.290 119.090 ;
        RECT 60.890 117.990 61.290 119.090 ;
        RECT 62.890 117.990 63.290 119.090 ;
        RECT 64.890 117.990 65.290 119.090 ;
        RECT 66.890 117.990 67.290 119.090 ;
        RECT 68.890 117.990 69.290 119.090 ;
        RECT 70.890 117.990 71.290 119.090 ;
        RECT 72.890 117.990 73.290 119.090 ;
        RECT 6.890 116.140 7.290 117.240 ;
        RECT 8.890 116.140 9.290 117.240 ;
        RECT 10.890 116.140 11.290 117.240 ;
        RECT 12.890 116.140 13.290 117.240 ;
        RECT 14.890 116.140 15.290 117.240 ;
        RECT 16.890 116.140 17.290 117.240 ;
        RECT 18.890 116.140 19.290 117.240 ;
        RECT 20.890 116.140 21.290 117.240 ;
        RECT 22.890 116.140 23.290 117.240 ;
        RECT 24.890 116.140 25.290 117.240 ;
        RECT 26.890 116.140 27.290 117.240 ;
        RECT 28.890 116.140 29.290 117.240 ;
        RECT 30.890 116.140 31.290 117.240 ;
        RECT 32.890 116.140 33.290 117.240 ;
        RECT 34.890 116.140 35.290 117.240 ;
        RECT 36.890 116.140 37.290 117.240 ;
        RECT 38.890 116.140 39.290 117.240 ;
        RECT 40.890 116.140 41.290 117.240 ;
        RECT 42.890 116.140 43.290 117.240 ;
        RECT 44.890 116.140 45.290 117.240 ;
        RECT 46.890 116.140 47.290 117.240 ;
        RECT 48.890 116.140 49.290 117.240 ;
        RECT 50.890 116.140 51.290 117.240 ;
        RECT 52.890 116.140 53.290 117.240 ;
        RECT 54.890 116.140 55.290 117.240 ;
        RECT 56.890 116.140 57.290 117.240 ;
        RECT 58.890 116.140 59.290 117.240 ;
        RECT 60.890 116.140 61.290 117.240 ;
        RECT 62.890 116.140 63.290 117.240 ;
        RECT 64.890 116.140 65.290 117.240 ;
        RECT 66.890 116.140 67.290 117.240 ;
        RECT 68.890 116.140 69.290 117.240 ;
        RECT 70.890 116.140 71.290 117.240 ;
        RECT 72.890 116.140 73.290 117.240 ;
        RECT 6.890 114.290 7.290 115.390 ;
        RECT 8.890 114.290 9.290 115.390 ;
        RECT 10.890 114.290 11.290 115.390 ;
        RECT 12.890 114.290 13.290 115.390 ;
        RECT 14.890 114.290 15.290 115.390 ;
        RECT 16.890 114.290 17.290 115.390 ;
        RECT 18.890 114.290 19.290 115.390 ;
        RECT 20.890 114.290 21.290 115.390 ;
        RECT 22.890 114.290 23.290 115.390 ;
        RECT 24.890 114.290 25.290 115.390 ;
        RECT 26.890 114.290 27.290 115.390 ;
        RECT 28.890 114.290 29.290 115.390 ;
        RECT 30.890 114.290 31.290 115.390 ;
        RECT 32.890 114.290 33.290 115.390 ;
        RECT 34.890 114.290 35.290 115.390 ;
        RECT 36.890 114.290 37.290 115.390 ;
        RECT 38.890 114.290 39.290 115.390 ;
        RECT 40.890 114.290 41.290 115.390 ;
        RECT 42.890 114.290 43.290 115.390 ;
        RECT 44.890 114.290 45.290 115.390 ;
        RECT 46.890 114.290 47.290 115.390 ;
        RECT 48.890 114.290 49.290 115.390 ;
        RECT 50.890 114.290 51.290 115.390 ;
        RECT 52.890 114.290 53.290 115.390 ;
        RECT 54.890 114.290 55.290 115.390 ;
        RECT 56.890 114.290 57.290 115.390 ;
        RECT 58.890 114.290 59.290 115.390 ;
        RECT 60.890 114.290 61.290 115.390 ;
        RECT 62.890 114.290 63.290 115.390 ;
        RECT 64.890 114.290 65.290 115.390 ;
        RECT 66.890 114.290 67.290 115.390 ;
        RECT 68.890 114.290 69.290 115.390 ;
        RECT 70.890 114.290 71.290 115.390 ;
        RECT 72.890 114.290 73.290 115.390 ;
        RECT 6.890 112.440 7.290 113.540 ;
        RECT 8.890 112.440 9.290 113.540 ;
        RECT 10.890 112.440 11.290 113.540 ;
        RECT 12.890 112.440 13.290 113.540 ;
        RECT 14.890 112.440 15.290 113.540 ;
        RECT 16.890 112.440 17.290 113.540 ;
        RECT 18.890 112.440 19.290 113.540 ;
        RECT 20.890 112.440 21.290 113.540 ;
        RECT 22.890 112.440 23.290 113.540 ;
        RECT 24.890 112.440 25.290 113.540 ;
        RECT 26.890 112.440 27.290 113.540 ;
        RECT 28.890 112.440 29.290 113.540 ;
        RECT 30.890 112.440 31.290 113.540 ;
        RECT 32.890 112.440 33.290 113.540 ;
        RECT 34.890 112.440 35.290 113.540 ;
        RECT 36.890 112.440 37.290 113.540 ;
        RECT 38.890 112.440 39.290 113.540 ;
        RECT 40.890 112.440 41.290 113.540 ;
        RECT 42.890 112.440 43.290 113.540 ;
        RECT 44.890 112.440 45.290 113.540 ;
        RECT 46.890 112.440 47.290 113.540 ;
        RECT 48.890 112.440 49.290 113.540 ;
        RECT 50.890 112.440 51.290 113.540 ;
        RECT 52.890 112.440 53.290 113.540 ;
        RECT 54.890 112.440 55.290 113.540 ;
        RECT 56.890 112.440 57.290 113.540 ;
        RECT 58.890 112.440 59.290 113.540 ;
        RECT 60.890 112.440 61.290 113.540 ;
        RECT 62.890 112.440 63.290 113.540 ;
        RECT 64.890 112.440 65.290 113.540 ;
        RECT 66.890 112.440 67.290 113.540 ;
        RECT 68.890 112.440 69.290 113.540 ;
        RECT 70.890 112.440 71.290 113.540 ;
        RECT 72.890 112.440 73.290 113.540 ;
        RECT 6.890 110.590 7.290 111.690 ;
        RECT 8.890 110.590 9.290 111.690 ;
        RECT 10.890 110.590 11.290 111.690 ;
        RECT 12.890 110.590 13.290 111.690 ;
        RECT 14.890 110.590 15.290 111.690 ;
        RECT 16.890 110.590 17.290 111.690 ;
        RECT 18.890 110.590 19.290 111.690 ;
        RECT 20.890 110.590 21.290 111.690 ;
        RECT 22.890 110.590 23.290 111.690 ;
        RECT 24.890 110.590 25.290 111.690 ;
        RECT 26.890 110.590 27.290 111.690 ;
        RECT 28.890 110.590 29.290 111.690 ;
        RECT 30.890 110.590 31.290 111.690 ;
        RECT 32.890 110.590 33.290 111.690 ;
        RECT 34.890 110.590 35.290 111.690 ;
        RECT 36.890 110.590 37.290 111.690 ;
        RECT 38.890 110.590 39.290 111.690 ;
        RECT 40.890 110.590 41.290 111.690 ;
        RECT 42.890 110.590 43.290 111.690 ;
        RECT 44.890 110.590 45.290 111.690 ;
        RECT 46.890 110.590 47.290 111.690 ;
        RECT 48.890 110.590 49.290 111.690 ;
        RECT 50.890 110.590 51.290 111.690 ;
        RECT 52.890 110.590 53.290 111.690 ;
        RECT 54.890 110.590 55.290 111.690 ;
        RECT 56.890 110.590 57.290 111.690 ;
        RECT 58.890 110.590 59.290 111.690 ;
        RECT 60.890 110.590 61.290 111.690 ;
        RECT 62.890 110.590 63.290 111.690 ;
        RECT 64.890 110.590 65.290 111.690 ;
        RECT 66.890 110.590 67.290 111.690 ;
        RECT 68.890 110.590 69.290 111.690 ;
        RECT 70.890 110.590 71.290 111.690 ;
        RECT 72.890 110.590 73.290 111.690 ;
        RECT 6.890 108.740 7.290 109.840 ;
        RECT 8.890 108.740 9.290 109.840 ;
        RECT 10.890 108.740 11.290 109.840 ;
        RECT 12.890 108.740 13.290 109.840 ;
        RECT 14.890 108.740 15.290 109.840 ;
        RECT 16.890 108.740 17.290 109.840 ;
        RECT 18.890 108.740 19.290 109.840 ;
        RECT 20.890 108.740 21.290 109.840 ;
        RECT 22.890 108.740 23.290 109.840 ;
        RECT 24.890 108.740 25.290 109.840 ;
        RECT 26.890 108.740 27.290 109.840 ;
        RECT 28.890 108.740 29.290 109.840 ;
        RECT 30.890 108.740 31.290 109.840 ;
        RECT 32.890 108.740 33.290 109.840 ;
        RECT 34.890 108.740 35.290 109.840 ;
        RECT 36.890 108.740 37.290 109.840 ;
        RECT 38.890 108.740 39.290 109.840 ;
        RECT 40.890 108.740 41.290 109.840 ;
        RECT 42.890 108.740 43.290 109.840 ;
        RECT 44.890 108.740 45.290 109.840 ;
        RECT 46.890 108.740 47.290 109.840 ;
        RECT 48.890 108.740 49.290 109.840 ;
        RECT 50.890 108.740 51.290 109.840 ;
        RECT 52.890 108.740 53.290 109.840 ;
        RECT 54.890 108.740 55.290 109.840 ;
        RECT 56.890 108.740 57.290 109.840 ;
        RECT 58.890 108.740 59.290 109.840 ;
        RECT 60.890 108.740 61.290 109.840 ;
        RECT 62.890 108.740 63.290 109.840 ;
        RECT 64.890 108.740 65.290 109.840 ;
        RECT 66.890 108.740 67.290 109.840 ;
        RECT 68.890 108.740 69.290 109.840 ;
        RECT 70.890 108.740 71.290 109.840 ;
        RECT 72.890 108.740 73.290 109.840 ;
        RECT 6.890 106.890 7.290 107.990 ;
        RECT 8.890 106.890 9.290 107.990 ;
        RECT 10.890 106.890 11.290 107.990 ;
        RECT 12.890 106.890 13.290 107.990 ;
        RECT 14.890 106.890 15.290 107.990 ;
        RECT 16.890 106.890 17.290 107.990 ;
        RECT 18.890 106.890 19.290 107.990 ;
        RECT 20.890 106.890 21.290 107.990 ;
        RECT 22.890 106.890 23.290 107.990 ;
        RECT 24.890 106.890 25.290 107.990 ;
        RECT 26.890 106.890 27.290 107.990 ;
        RECT 28.890 106.890 29.290 107.990 ;
        RECT 30.890 106.890 31.290 107.990 ;
        RECT 32.890 106.890 33.290 107.990 ;
        RECT 34.890 106.890 35.290 107.990 ;
        RECT 36.890 106.890 37.290 107.990 ;
        RECT 38.890 106.890 39.290 107.990 ;
        RECT 40.890 106.890 41.290 107.990 ;
        RECT 42.890 106.890 43.290 107.990 ;
        RECT 44.890 106.890 45.290 107.990 ;
        RECT 46.890 106.890 47.290 107.990 ;
        RECT 48.890 106.890 49.290 107.990 ;
        RECT 50.890 106.890 51.290 107.990 ;
        RECT 52.890 106.890 53.290 107.990 ;
        RECT 54.890 106.890 55.290 107.990 ;
        RECT 56.890 106.890 57.290 107.990 ;
        RECT 58.890 106.890 59.290 107.990 ;
        RECT 60.890 106.890 61.290 107.990 ;
        RECT 62.890 106.890 63.290 107.990 ;
        RECT 64.890 106.890 65.290 107.990 ;
        RECT 66.890 106.890 67.290 107.990 ;
        RECT 68.890 106.890 69.290 107.990 ;
        RECT 70.890 106.890 71.290 107.990 ;
        RECT 72.890 106.890 73.290 107.990 ;
        RECT 6.890 105.040 7.290 106.140 ;
        RECT 8.890 105.040 9.290 106.140 ;
        RECT 10.890 105.040 11.290 106.140 ;
        RECT 12.890 105.040 13.290 106.140 ;
        RECT 14.890 105.040 15.290 106.140 ;
        RECT 16.890 105.040 17.290 106.140 ;
        RECT 18.890 105.040 19.290 106.140 ;
        RECT 20.890 105.040 21.290 106.140 ;
        RECT 22.890 105.040 23.290 106.140 ;
        RECT 24.890 105.040 25.290 106.140 ;
        RECT 26.890 105.040 27.290 106.140 ;
        RECT 28.890 105.040 29.290 106.140 ;
        RECT 30.890 105.040 31.290 106.140 ;
        RECT 32.890 105.040 33.290 106.140 ;
        RECT 34.890 105.040 35.290 106.140 ;
        RECT 36.890 105.040 37.290 106.140 ;
        RECT 38.890 105.040 39.290 106.140 ;
        RECT 40.890 105.040 41.290 106.140 ;
        RECT 42.890 105.040 43.290 106.140 ;
        RECT 44.890 105.040 45.290 106.140 ;
        RECT 46.890 105.040 47.290 106.140 ;
        RECT 48.890 105.040 49.290 106.140 ;
        RECT 50.890 105.040 51.290 106.140 ;
        RECT 52.890 105.040 53.290 106.140 ;
        RECT 54.890 105.040 55.290 106.140 ;
        RECT 56.890 105.040 57.290 106.140 ;
        RECT 58.890 105.040 59.290 106.140 ;
        RECT 60.890 105.040 61.290 106.140 ;
        RECT 62.890 105.040 63.290 106.140 ;
        RECT 64.890 105.040 65.290 106.140 ;
        RECT 66.890 105.040 67.290 106.140 ;
        RECT 68.890 105.040 69.290 106.140 ;
        RECT 70.890 105.040 71.290 106.140 ;
        RECT 72.890 105.040 73.290 106.140 ;
        RECT 6.890 103.190 7.290 104.290 ;
        RECT 8.890 103.190 9.290 104.290 ;
        RECT 10.890 103.190 11.290 104.290 ;
        RECT 12.890 103.190 13.290 104.290 ;
        RECT 14.890 103.190 15.290 104.290 ;
        RECT 16.890 103.190 17.290 104.290 ;
        RECT 18.890 103.190 19.290 104.290 ;
        RECT 20.890 103.190 21.290 104.290 ;
        RECT 22.890 103.190 23.290 104.290 ;
        RECT 24.890 103.190 25.290 104.290 ;
        RECT 26.890 103.190 27.290 104.290 ;
        RECT 28.890 103.190 29.290 104.290 ;
        RECT 30.890 103.190 31.290 104.290 ;
        RECT 32.890 103.190 33.290 104.290 ;
        RECT 34.890 103.190 35.290 104.290 ;
        RECT 36.890 103.190 37.290 104.290 ;
        RECT 38.890 103.190 39.290 104.290 ;
        RECT 40.890 103.190 41.290 104.290 ;
        RECT 42.890 103.190 43.290 104.290 ;
        RECT 44.890 103.190 45.290 104.290 ;
        RECT 46.890 103.190 47.290 104.290 ;
        RECT 48.890 103.190 49.290 104.290 ;
        RECT 50.890 103.190 51.290 104.290 ;
        RECT 52.890 103.190 53.290 104.290 ;
        RECT 54.890 103.190 55.290 104.290 ;
        RECT 56.890 103.190 57.290 104.290 ;
        RECT 58.890 103.190 59.290 104.290 ;
        RECT 60.890 103.190 61.290 104.290 ;
        RECT 62.890 103.190 63.290 104.290 ;
        RECT 64.890 103.190 65.290 104.290 ;
        RECT 66.890 103.190 67.290 104.290 ;
        RECT 68.890 103.190 69.290 104.290 ;
        RECT 70.890 103.190 71.290 104.290 ;
        RECT 72.890 103.190 73.290 104.290 ;
        RECT 6.890 101.340 7.290 102.440 ;
        RECT 8.890 101.340 9.290 102.440 ;
        RECT 10.890 101.340 11.290 102.440 ;
        RECT 12.890 101.340 13.290 102.440 ;
        RECT 14.890 101.340 15.290 102.440 ;
        RECT 16.890 101.340 17.290 102.440 ;
        RECT 18.890 101.340 19.290 102.440 ;
        RECT 20.890 101.340 21.290 102.440 ;
        RECT 22.890 101.340 23.290 102.440 ;
        RECT 24.890 101.340 25.290 102.440 ;
        RECT 26.890 101.340 27.290 102.440 ;
        RECT 28.890 101.340 29.290 102.440 ;
        RECT 30.890 101.340 31.290 102.440 ;
        RECT 32.890 101.340 33.290 102.440 ;
        RECT 34.890 101.340 35.290 102.440 ;
        RECT 36.890 101.340 37.290 102.440 ;
        RECT 38.890 101.340 39.290 102.440 ;
        RECT 40.890 101.340 41.290 102.440 ;
        RECT 42.890 101.340 43.290 102.440 ;
        RECT 44.890 101.340 45.290 102.440 ;
        RECT 46.890 101.340 47.290 102.440 ;
        RECT 48.890 101.340 49.290 102.440 ;
        RECT 50.890 101.340 51.290 102.440 ;
        RECT 52.890 101.340 53.290 102.440 ;
        RECT 54.890 101.340 55.290 102.440 ;
        RECT 56.890 101.340 57.290 102.440 ;
        RECT 58.890 101.340 59.290 102.440 ;
        RECT 60.890 101.340 61.290 102.440 ;
        RECT 62.890 101.340 63.290 102.440 ;
        RECT 64.890 101.340 65.290 102.440 ;
        RECT 66.890 101.340 67.290 102.440 ;
        RECT 68.890 101.340 69.290 102.440 ;
        RECT 70.890 101.340 71.290 102.440 ;
        RECT 72.890 101.340 73.290 102.440 ;
        RECT 6.890 99.490 7.290 100.590 ;
        RECT 8.890 99.490 9.290 100.590 ;
        RECT 10.890 99.490 11.290 100.590 ;
        RECT 12.890 99.490 13.290 100.590 ;
        RECT 14.890 99.490 15.290 100.590 ;
        RECT 16.890 99.490 17.290 100.590 ;
        RECT 18.890 99.490 19.290 100.590 ;
        RECT 20.890 99.490 21.290 100.590 ;
        RECT 22.890 99.490 23.290 100.590 ;
        RECT 24.890 99.490 25.290 100.590 ;
        RECT 26.890 99.490 27.290 100.590 ;
        RECT 28.890 99.490 29.290 100.590 ;
        RECT 30.890 99.490 31.290 100.590 ;
        RECT 32.890 99.490 33.290 100.590 ;
        RECT 34.890 99.490 35.290 100.590 ;
        RECT 36.890 99.490 37.290 100.590 ;
        RECT 38.890 99.490 39.290 100.590 ;
        RECT 40.890 99.490 41.290 100.590 ;
        RECT 42.890 99.490 43.290 100.590 ;
        RECT 44.890 99.490 45.290 100.590 ;
        RECT 46.890 99.490 47.290 100.590 ;
        RECT 48.890 99.490 49.290 100.590 ;
        RECT 50.890 99.490 51.290 100.590 ;
        RECT 52.890 99.490 53.290 100.590 ;
        RECT 54.890 99.490 55.290 100.590 ;
        RECT 56.890 99.490 57.290 100.590 ;
        RECT 58.890 99.490 59.290 100.590 ;
        RECT 60.890 99.490 61.290 100.590 ;
        RECT 62.890 99.490 63.290 100.590 ;
        RECT 64.890 99.490 65.290 100.590 ;
        RECT 66.890 99.490 67.290 100.590 ;
        RECT 68.890 99.490 69.290 100.590 ;
        RECT 70.890 99.490 71.290 100.590 ;
        RECT 72.890 99.490 73.290 100.590 ;
        RECT 6.890 97.640 7.290 98.740 ;
        RECT 8.890 97.640 9.290 98.740 ;
        RECT 10.890 97.640 11.290 98.740 ;
        RECT 12.890 97.640 13.290 98.740 ;
        RECT 14.890 97.640 15.290 98.740 ;
        RECT 16.890 97.640 17.290 98.740 ;
        RECT 18.890 97.640 19.290 98.740 ;
        RECT 20.890 97.640 21.290 98.740 ;
        RECT 22.890 97.640 23.290 98.740 ;
        RECT 24.890 97.640 25.290 98.740 ;
        RECT 26.890 97.640 27.290 98.740 ;
        RECT 28.890 97.640 29.290 98.740 ;
        RECT 30.890 97.640 31.290 98.740 ;
        RECT 32.890 97.640 33.290 98.740 ;
        RECT 34.890 97.640 35.290 98.740 ;
        RECT 36.890 97.640 37.290 98.740 ;
        RECT 38.890 97.640 39.290 98.740 ;
        RECT 40.890 97.640 41.290 98.740 ;
        RECT 42.890 97.640 43.290 98.740 ;
        RECT 44.890 97.640 45.290 98.740 ;
        RECT 46.890 97.640 47.290 98.740 ;
        RECT 48.890 97.640 49.290 98.740 ;
        RECT 50.890 97.640 51.290 98.740 ;
        RECT 52.890 97.640 53.290 98.740 ;
        RECT 54.890 97.640 55.290 98.740 ;
        RECT 56.890 97.640 57.290 98.740 ;
        RECT 58.890 97.640 59.290 98.740 ;
        RECT 60.890 97.640 61.290 98.740 ;
        RECT 62.890 97.640 63.290 98.740 ;
        RECT 64.890 97.640 65.290 98.740 ;
        RECT 66.890 97.640 67.290 98.740 ;
        RECT 68.890 97.640 69.290 98.740 ;
        RECT 70.890 97.640 71.290 98.740 ;
        RECT 72.890 97.640 73.290 98.740 ;
        RECT 6.890 95.790 7.290 96.890 ;
        RECT 8.890 95.790 9.290 96.890 ;
        RECT 10.890 95.790 11.290 96.890 ;
        RECT 12.890 95.790 13.290 96.890 ;
        RECT 14.890 95.790 15.290 96.890 ;
        RECT 16.890 95.790 17.290 96.890 ;
        RECT 18.890 95.790 19.290 96.890 ;
        RECT 20.890 95.790 21.290 96.890 ;
        RECT 22.890 95.790 23.290 96.890 ;
        RECT 24.890 95.790 25.290 96.890 ;
        RECT 26.890 95.790 27.290 96.890 ;
        RECT 28.890 95.790 29.290 96.890 ;
        RECT 30.890 95.790 31.290 96.890 ;
        RECT 32.890 95.790 33.290 96.890 ;
        RECT 34.890 95.790 35.290 96.890 ;
        RECT 36.890 95.790 37.290 96.890 ;
        RECT 38.890 95.790 39.290 96.890 ;
        RECT 40.890 95.790 41.290 96.890 ;
        RECT 42.890 95.790 43.290 96.890 ;
        RECT 44.890 95.790 45.290 96.890 ;
        RECT 46.890 95.790 47.290 96.890 ;
        RECT 48.890 95.790 49.290 96.890 ;
        RECT 50.890 95.790 51.290 96.890 ;
        RECT 52.890 95.790 53.290 96.890 ;
        RECT 54.890 95.790 55.290 96.890 ;
        RECT 56.890 95.790 57.290 96.890 ;
        RECT 58.890 95.790 59.290 96.890 ;
        RECT 60.890 95.790 61.290 96.890 ;
        RECT 62.890 95.790 63.290 96.890 ;
        RECT 64.890 95.790 65.290 96.890 ;
        RECT 66.890 95.790 67.290 96.890 ;
        RECT 68.890 95.790 69.290 96.890 ;
        RECT 70.890 95.790 71.290 96.890 ;
        RECT 72.890 95.790 73.290 96.890 ;
        RECT 6.890 93.940 7.290 95.040 ;
        RECT 8.890 93.940 9.290 95.040 ;
        RECT 10.890 93.940 11.290 95.040 ;
        RECT 12.890 93.940 13.290 95.040 ;
        RECT 14.890 93.940 15.290 95.040 ;
        RECT 16.890 93.940 17.290 95.040 ;
        RECT 18.890 93.940 19.290 95.040 ;
        RECT 20.890 93.940 21.290 95.040 ;
        RECT 22.890 93.940 23.290 95.040 ;
        RECT 24.890 93.940 25.290 95.040 ;
        RECT 26.890 93.940 27.290 95.040 ;
        RECT 28.890 93.940 29.290 95.040 ;
        RECT 30.890 93.940 31.290 95.040 ;
        RECT 32.890 93.940 33.290 95.040 ;
        RECT 34.890 93.940 35.290 95.040 ;
        RECT 36.890 93.940 37.290 95.040 ;
        RECT 38.890 93.940 39.290 95.040 ;
        RECT 40.890 93.940 41.290 95.040 ;
        RECT 42.890 93.940 43.290 95.040 ;
        RECT 44.890 93.940 45.290 95.040 ;
        RECT 46.890 93.940 47.290 95.040 ;
        RECT 48.890 93.940 49.290 95.040 ;
        RECT 50.890 93.940 51.290 95.040 ;
        RECT 52.890 93.940 53.290 95.040 ;
        RECT 54.890 93.940 55.290 95.040 ;
        RECT 56.890 93.940 57.290 95.040 ;
        RECT 58.890 93.940 59.290 95.040 ;
        RECT 60.890 93.940 61.290 95.040 ;
        RECT 62.890 93.940 63.290 95.040 ;
        RECT 64.890 93.940 65.290 95.040 ;
        RECT 66.890 93.940 67.290 95.040 ;
        RECT 68.890 93.940 69.290 95.040 ;
        RECT 70.890 93.940 71.290 95.040 ;
        RECT 72.890 93.940 73.290 95.040 ;
        RECT 6.890 92.090 7.290 93.190 ;
        RECT 8.890 92.090 9.290 93.190 ;
        RECT 10.890 92.090 11.290 93.190 ;
        RECT 12.890 92.090 13.290 93.190 ;
        RECT 14.890 92.090 15.290 93.190 ;
        RECT 16.890 92.090 17.290 93.190 ;
        RECT 18.890 92.090 19.290 93.190 ;
        RECT 20.890 92.090 21.290 93.190 ;
        RECT 22.890 92.090 23.290 93.190 ;
        RECT 24.890 92.090 25.290 93.190 ;
        RECT 26.890 92.090 27.290 93.190 ;
        RECT 28.890 92.090 29.290 93.190 ;
        RECT 30.890 92.090 31.290 93.190 ;
        RECT 32.890 92.090 33.290 93.190 ;
        RECT 34.890 92.090 35.290 93.190 ;
        RECT 36.890 92.090 37.290 93.190 ;
        RECT 38.890 92.090 39.290 93.190 ;
        RECT 40.890 92.090 41.290 93.190 ;
        RECT 42.890 92.090 43.290 93.190 ;
        RECT 44.890 92.090 45.290 93.190 ;
        RECT 46.890 92.090 47.290 93.190 ;
        RECT 48.890 92.090 49.290 93.190 ;
        RECT 50.890 92.090 51.290 93.190 ;
        RECT 52.890 92.090 53.290 93.190 ;
        RECT 54.890 92.090 55.290 93.190 ;
        RECT 56.890 92.090 57.290 93.190 ;
        RECT 58.890 92.090 59.290 93.190 ;
        RECT 60.890 92.090 61.290 93.190 ;
        RECT 62.890 92.090 63.290 93.190 ;
        RECT 64.890 92.090 65.290 93.190 ;
        RECT 66.890 92.090 67.290 93.190 ;
        RECT 68.890 92.090 69.290 93.190 ;
        RECT 70.890 92.090 71.290 93.190 ;
        RECT 72.890 92.090 73.290 93.190 ;
        RECT 6.890 90.240 7.290 91.340 ;
        RECT 8.890 90.240 9.290 91.340 ;
        RECT 10.890 90.240 11.290 91.340 ;
        RECT 12.890 90.240 13.290 91.340 ;
        RECT 14.890 90.240 15.290 91.340 ;
        RECT 16.890 90.240 17.290 91.340 ;
        RECT 18.890 90.240 19.290 91.340 ;
        RECT 20.890 90.240 21.290 91.340 ;
        RECT 22.890 90.240 23.290 91.340 ;
        RECT 24.890 90.240 25.290 91.340 ;
        RECT 26.890 90.240 27.290 91.340 ;
        RECT 28.890 90.240 29.290 91.340 ;
        RECT 30.890 90.240 31.290 91.340 ;
        RECT 32.890 90.240 33.290 91.340 ;
        RECT 34.890 90.240 35.290 91.340 ;
        RECT 36.890 90.240 37.290 91.340 ;
        RECT 38.890 90.240 39.290 91.340 ;
        RECT 40.890 90.240 41.290 91.340 ;
        RECT 42.890 90.240 43.290 91.340 ;
        RECT 44.890 90.240 45.290 91.340 ;
        RECT 46.890 90.240 47.290 91.340 ;
        RECT 48.890 90.240 49.290 91.340 ;
        RECT 50.890 90.240 51.290 91.340 ;
        RECT 52.890 90.240 53.290 91.340 ;
        RECT 54.890 90.240 55.290 91.340 ;
        RECT 56.890 90.240 57.290 91.340 ;
        RECT 58.890 90.240 59.290 91.340 ;
        RECT 60.890 90.240 61.290 91.340 ;
        RECT 62.890 90.240 63.290 91.340 ;
        RECT 64.890 90.240 65.290 91.340 ;
        RECT 66.890 90.240 67.290 91.340 ;
        RECT 68.890 90.240 69.290 91.340 ;
        RECT 70.890 90.240 71.290 91.340 ;
        RECT 72.890 90.240 73.290 91.340 ;
        RECT 6.890 88.390 7.290 89.490 ;
        RECT 8.890 88.390 9.290 89.490 ;
        RECT 10.890 88.390 11.290 89.490 ;
        RECT 12.890 88.390 13.290 89.490 ;
        RECT 14.890 88.390 15.290 89.490 ;
        RECT 16.890 88.390 17.290 89.490 ;
        RECT 18.890 88.390 19.290 89.490 ;
        RECT 20.890 88.390 21.290 89.490 ;
        RECT 22.890 88.390 23.290 89.490 ;
        RECT 24.890 88.390 25.290 89.490 ;
        RECT 26.890 88.390 27.290 89.490 ;
        RECT 28.890 88.390 29.290 89.490 ;
        RECT 30.890 88.390 31.290 89.490 ;
        RECT 32.890 88.390 33.290 89.490 ;
        RECT 34.890 88.390 35.290 89.490 ;
        RECT 36.890 88.390 37.290 89.490 ;
        RECT 38.890 88.390 39.290 89.490 ;
        RECT 40.890 88.390 41.290 89.490 ;
        RECT 42.890 88.390 43.290 89.490 ;
        RECT 44.890 88.390 45.290 89.490 ;
        RECT 46.890 88.390 47.290 89.490 ;
        RECT 48.890 88.390 49.290 89.490 ;
        RECT 50.890 88.390 51.290 89.490 ;
        RECT 52.890 88.390 53.290 89.490 ;
        RECT 54.890 88.390 55.290 89.490 ;
        RECT 56.890 88.390 57.290 89.490 ;
        RECT 58.890 88.390 59.290 89.490 ;
        RECT 60.890 88.390 61.290 89.490 ;
        RECT 62.890 88.390 63.290 89.490 ;
        RECT 64.890 88.390 65.290 89.490 ;
        RECT 66.890 88.390 67.290 89.490 ;
        RECT 68.890 88.390 69.290 89.490 ;
        RECT 70.890 88.390 71.290 89.490 ;
        RECT 72.890 88.390 73.290 89.490 ;
        RECT 6.890 86.540 7.290 87.640 ;
        RECT 8.890 86.540 9.290 87.640 ;
        RECT 10.890 86.540 11.290 87.640 ;
        RECT 12.890 86.540 13.290 87.640 ;
        RECT 14.890 86.540 15.290 87.640 ;
        RECT 16.890 86.540 17.290 87.640 ;
        RECT 18.890 86.540 19.290 87.640 ;
        RECT 20.890 86.540 21.290 87.640 ;
        RECT 22.890 86.540 23.290 87.640 ;
        RECT 24.890 86.540 25.290 87.640 ;
        RECT 26.890 86.540 27.290 87.640 ;
        RECT 28.890 86.540 29.290 87.640 ;
        RECT 30.890 86.540 31.290 87.640 ;
        RECT 32.890 86.540 33.290 87.640 ;
        RECT 34.890 86.540 35.290 87.640 ;
        RECT 36.890 86.540 37.290 87.640 ;
        RECT 38.890 86.540 39.290 87.640 ;
        RECT 40.890 86.540 41.290 87.640 ;
        RECT 42.890 86.540 43.290 87.640 ;
        RECT 44.890 86.540 45.290 87.640 ;
        RECT 46.890 86.540 47.290 87.640 ;
        RECT 48.890 86.540 49.290 87.640 ;
        RECT 50.890 86.540 51.290 87.640 ;
        RECT 52.890 86.540 53.290 87.640 ;
        RECT 54.890 86.540 55.290 87.640 ;
        RECT 56.890 86.540 57.290 87.640 ;
        RECT 58.890 86.540 59.290 87.640 ;
        RECT 60.890 86.540 61.290 87.640 ;
        RECT 62.890 86.540 63.290 87.640 ;
        RECT 64.890 86.540 65.290 87.640 ;
        RECT 66.890 86.540 67.290 87.640 ;
        RECT 68.890 86.540 69.290 87.640 ;
        RECT 70.890 86.540 71.290 87.640 ;
        RECT 72.890 86.540 73.290 87.640 ;
        RECT 6.890 84.690 7.290 85.790 ;
        RECT 8.890 84.690 9.290 85.790 ;
        RECT 10.890 84.690 11.290 85.790 ;
        RECT 12.890 84.690 13.290 85.790 ;
        RECT 14.890 84.690 15.290 85.790 ;
        RECT 16.890 84.690 17.290 85.790 ;
        RECT 18.890 84.690 19.290 85.790 ;
        RECT 20.890 84.690 21.290 85.790 ;
        RECT 22.890 84.690 23.290 85.790 ;
        RECT 24.890 84.690 25.290 85.790 ;
        RECT 26.890 84.690 27.290 85.790 ;
        RECT 28.890 84.690 29.290 85.790 ;
        RECT 30.890 84.690 31.290 85.790 ;
        RECT 32.890 84.690 33.290 85.790 ;
        RECT 34.890 84.690 35.290 85.790 ;
        RECT 36.890 84.690 37.290 85.790 ;
        RECT 38.890 84.690 39.290 85.790 ;
        RECT 40.890 84.690 41.290 85.790 ;
        RECT 42.890 84.690 43.290 85.790 ;
        RECT 44.890 84.690 45.290 85.790 ;
        RECT 46.890 84.690 47.290 85.790 ;
        RECT 48.890 84.690 49.290 85.790 ;
        RECT 50.890 84.690 51.290 85.790 ;
        RECT 52.890 84.690 53.290 85.790 ;
        RECT 54.890 84.690 55.290 85.790 ;
        RECT 56.890 84.690 57.290 85.790 ;
        RECT 58.890 84.690 59.290 85.790 ;
        RECT 60.890 84.690 61.290 85.790 ;
        RECT 62.890 84.690 63.290 85.790 ;
        RECT 64.890 84.690 65.290 85.790 ;
        RECT 66.890 84.690 67.290 85.790 ;
        RECT 68.890 84.690 69.290 85.790 ;
        RECT 70.890 84.690 71.290 85.790 ;
        RECT 72.890 84.690 73.290 85.790 ;
        RECT 6.890 82.840 7.290 83.940 ;
        RECT 8.890 82.840 9.290 83.940 ;
        RECT 10.890 82.840 11.290 83.940 ;
        RECT 12.890 82.840 13.290 83.940 ;
        RECT 14.890 82.840 15.290 83.940 ;
        RECT 16.890 82.840 17.290 83.940 ;
        RECT 18.890 82.840 19.290 83.940 ;
        RECT 20.890 82.840 21.290 83.940 ;
        RECT 22.890 82.840 23.290 83.940 ;
        RECT 24.890 82.840 25.290 83.940 ;
        RECT 26.890 82.840 27.290 83.940 ;
        RECT 28.890 82.840 29.290 83.940 ;
        RECT 30.890 82.840 31.290 83.940 ;
        RECT 32.890 82.840 33.290 83.940 ;
        RECT 34.890 82.840 35.290 83.940 ;
        RECT 36.890 82.840 37.290 83.940 ;
        RECT 38.890 82.840 39.290 83.940 ;
        RECT 40.890 82.840 41.290 83.940 ;
        RECT 42.890 82.840 43.290 83.940 ;
        RECT 44.890 82.840 45.290 83.940 ;
        RECT 46.890 82.840 47.290 83.940 ;
        RECT 48.890 82.840 49.290 83.940 ;
        RECT 50.890 82.840 51.290 83.940 ;
        RECT 52.890 82.840 53.290 83.940 ;
        RECT 54.890 82.840 55.290 83.940 ;
        RECT 56.890 82.840 57.290 83.940 ;
        RECT 58.890 82.840 59.290 83.940 ;
        RECT 60.890 82.840 61.290 83.940 ;
        RECT 62.890 82.840 63.290 83.940 ;
        RECT 64.890 82.840 65.290 83.940 ;
        RECT 66.890 82.840 67.290 83.940 ;
        RECT 68.890 82.840 69.290 83.940 ;
        RECT 70.890 82.840 71.290 83.940 ;
        RECT 72.890 82.840 73.290 83.940 ;
        RECT 6.890 80.990 7.290 82.090 ;
        RECT 8.890 80.990 9.290 82.090 ;
        RECT 10.890 80.990 11.290 82.090 ;
        RECT 12.890 80.990 13.290 82.090 ;
        RECT 14.890 80.990 15.290 82.090 ;
        RECT 16.890 80.990 17.290 82.090 ;
        RECT 18.890 80.990 19.290 82.090 ;
        RECT 20.890 80.990 21.290 82.090 ;
        RECT 22.890 80.990 23.290 82.090 ;
        RECT 24.890 80.990 25.290 82.090 ;
        RECT 26.890 80.990 27.290 82.090 ;
        RECT 28.890 80.990 29.290 82.090 ;
        RECT 30.890 80.990 31.290 82.090 ;
        RECT 32.890 80.990 33.290 82.090 ;
        RECT 34.890 80.990 35.290 82.090 ;
        RECT 36.890 80.990 37.290 82.090 ;
        RECT 38.890 80.990 39.290 82.090 ;
        RECT 40.890 80.990 41.290 82.090 ;
        RECT 42.890 80.990 43.290 82.090 ;
        RECT 44.890 80.990 45.290 82.090 ;
        RECT 46.890 80.990 47.290 82.090 ;
        RECT 48.890 80.990 49.290 82.090 ;
        RECT 50.890 80.990 51.290 82.090 ;
        RECT 52.890 80.990 53.290 82.090 ;
        RECT 54.890 80.990 55.290 82.090 ;
        RECT 56.890 80.990 57.290 82.090 ;
        RECT 58.890 80.990 59.290 82.090 ;
        RECT 60.890 80.990 61.290 82.090 ;
        RECT 62.890 80.990 63.290 82.090 ;
        RECT 64.890 80.990 65.290 82.090 ;
        RECT 66.890 80.990 67.290 82.090 ;
        RECT 68.890 80.990 69.290 82.090 ;
        RECT 70.890 80.990 71.290 82.090 ;
        RECT 72.890 80.990 73.290 82.090 ;
        RECT 6.890 79.140 7.290 80.240 ;
        RECT 8.890 79.140 9.290 80.240 ;
        RECT 10.890 79.140 11.290 80.240 ;
        RECT 12.890 79.140 13.290 80.240 ;
        RECT 14.890 79.140 15.290 80.240 ;
        RECT 16.890 79.140 17.290 80.240 ;
        RECT 18.890 79.140 19.290 80.240 ;
        RECT 20.890 79.140 21.290 80.240 ;
        RECT 22.890 79.140 23.290 80.240 ;
        RECT 24.890 79.140 25.290 80.240 ;
        RECT 26.890 79.140 27.290 80.240 ;
        RECT 28.890 79.140 29.290 80.240 ;
        RECT 30.890 79.140 31.290 80.240 ;
        RECT 32.890 79.140 33.290 80.240 ;
        RECT 34.890 79.140 35.290 80.240 ;
        RECT 36.890 79.140 37.290 80.240 ;
        RECT 38.890 79.140 39.290 80.240 ;
        RECT 40.890 79.140 41.290 80.240 ;
        RECT 42.890 79.140 43.290 80.240 ;
        RECT 44.890 79.140 45.290 80.240 ;
        RECT 46.890 79.140 47.290 80.240 ;
        RECT 48.890 79.140 49.290 80.240 ;
        RECT 50.890 79.140 51.290 80.240 ;
        RECT 52.890 79.140 53.290 80.240 ;
        RECT 54.890 79.140 55.290 80.240 ;
        RECT 56.890 79.140 57.290 80.240 ;
        RECT 58.890 79.140 59.290 80.240 ;
        RECT 60.890 79.140 61.290 80.240 ;
        RECT 62.890 79.140 63.290 80.240 ;
        RECT 64.890 79.140 65.290 80.240 ;
        RECT 66.890 79.140 67.290 80.240 ;
        RECT 68.890 79.140 69.290 80.240 ;
        RECT 70.890 79.140 71.290 80.240 ;
        RECT 72.890 79.140 73.290 80.240 ;
        RECT 6.890 77.290 7.290 78.390 ;
        RECT 8.890 77.290 9.290 78.390 ;
        RECT 10.890 77.290 11.290 78.390 ;
        RECT 12.890 77.290 13.290 78.390 ;
        RECT 14.890 77.290 15.290 78.390 ;
        RECT 16.890 77.290 17.290 78.390 ;
        RECT 18.890 77.290 19.290 78.390 ;
        RECT 20.890 77.290 21.290 78.390 ;
        RECT 22.890 77.290 23.290 78.390 ;
        RECT 24.890 77.290 25.290 78.390 ;
        RECT 26.890 77.290 27.290 78.390 ;
        RECT 28.890 77.290 29.290 78.390 ;
        RECT 30.890 77.290 31.290 78.390 ;
        RECT 32.890 77.290 33.290 78.390 ;
        RECT 34.890 77.290 35.290 78.390 ;
        RECT 36.890 77.290 37.290 78.390 ;
        RECT 38.890 77.290 39.290 78.390 ;
        RECT 40.890 77.290 41.290 78.390 ;
        RECT 42.890 77.290 43.290 78.390 ;
        RECT 44.890 77.290 45.290 78.390 ;
        RECT 46.890 77.290 47.290 78.390 ;
        RECT 48.890 77.290 49.290 78.390 ;
        RECT 50.890 77.290 51.290 78.390 ;
        RECT 52.890 77.290 53.290 78.390 ;
        RECT 54.890 77.290 55.290 78.390 ;
        RECT 56.890 77.290 57.290 78.390 ;
        RECT 58.890 77.290 59.290 78.390 ;
        RECT 60.890 77.290 61.290 78.390 ;
        RECT 62.890 77.290 63.290 78.390 ;
        RECT 64.890 77.290 65.290 78.390 ;
        RECT 66.890 77.290 67.290 78.390 ;
        RECT 68.890 77.290 69.290 78.390 ;
        RECT 70.890 77.290 71.290 78.390 ;
        RECT 72.890 77.290 73.290 78.390 ;
        RECT 6.890 75.440 7.290 76.540 ;
        RECT 8.890 75.440 9.290 76.540 ;
        RECT 10.890 75.440 11.290 76.540 ;
        RECT 12.890 75.440 13.290 76.540 ;
        RECT 14.890 75.440 15.290 76.540 ;
        RECT 16.890 75.440 17.290 76.540 ;
        RECT 18.890 75.440 19.290 76.540 ;
        RECT 20.890 75.440 21.290 76.540 ;
        RECT 22.890 75.440 23.290 76.540 ;
        RECT 24.890 75.440 25.290 76.540 ;
        RECT 26.890 75.440 27.290 76.540 ;
        RECT 28.890 75.440 29.290 76.540 ;
        RECT 30.890 75.440 31.290 76.540 ;
        RECT 32.890 75.440 33.290 76.540 ;
        RECT 34.890 75.440 35.290 76.540 ;
        RECT 36.890 75.440 37.290 76.540 ;
        RECT 38.890 75.440 39.290 76.540 ;
        RECT 40.890 75.440 41.290 76.540 ;
        RECT 42.890 75.440 43.290 76.540 ;
        RECT 44.890 75.440 45.290 76.540 ;
        RECT 46.890 75.440 47.290 76.540 ;
        RECT 48.890 75.440 49.290 76.540 ;
        RECT 50.890 75.440 51.290 76.540 ;
        RECT 52.890 75.440 53.290 76.540 ;
        RECT 54.890 75.440 55.290 76.540 ;
        RECT 56.890 75.440 57.290 76.540 ;
        RECT 58.890 75.440 59.290 76.540 ;
        RECT 60.890 75.440 61.290 76.540 ;
        RECT 62.890 75.440 63.290 76.540 ;
        RECT 64.890 75.440 65.290 76.540 ;
        RECT 66.890 75.440 67.290 76.540 ;
        RECT 68.890 75.440 69.290 76.540 ;
        RECT 70.890 75.440 71.290 76.540 ;
        RECT 72.890 75.440 73.290 76.540 ;
        RECT 6.890 73.590 7.290 74.690 ;
        RECT 8.890 73.590 9.290 74.690 ;
        RECT 10.890 73.590 11.290 74.690 ;
        RECT 12.890 73.590 13.290 74.690 ;
        RECT 14.890 73.590 15.290 74.690 ;
        RECT 16.890 73.590 17.290 74.690 ;
        RECT 18.890 73.590 19.290 74.690 ;
        RECT 20.890 73.590 21.290 74.690 ;
        RECT 22.890 73.590 23.290 74.690 ;
        RECT 24.890 73.590 25.290 74.690 ;
        RECT 26.890 73.590 27.290 74.690 ;
        RECT 28.890 73.590 29.290 74.690 ;
        RECT 30.890 73.590 31.290 74.690 ;
        RECT 32.890 73.590 33.290 74.690 ;
        RECT 34.890 73.590 35.290 74.690 ;
        RECT 36.890 73.590 37.290 74.690 ;
        RECT 38.890 73.590 39.290 74.690 ;
        RECT 40.890 73.590 41.290 74.690 ;
        RECT 42.890 73.590 43.290 74.690 ;
        RECT 44.890 73.590 45.290 74.690 ;
        RECT 46.890 73.590 47.290 74.690 ;
        RECT 48.890 73.590 49.290 74.690 ;
        RECT 50.890 73.590 51.290 74.690 ;
        RECT 52.890 73.590 53.290 74.690 ;
        RECT 54.890 73.590 55.290 74.690 ;
        RECT 56.890 73.590 57.290 74.690 ;
        RECT 58.890 73.590 59.290 74.690 ;
        RECT 60.890 73.590 61.290 74.690 ;
        RECT 62.890 73.590 63.290 74.690 ;
        RECT 64.890 73.590 65.290 74.690 ;
        RECT 66.890 73.590 67.290 74.690 ;
        RECT 68.890 73.590 69.290 74.690 ;
        RECT 70.890 73.590 71.290 74.690 ;
        RECT 72.890 73.590 73.290 74.690 ;
        RECT 6.890 71.740 7.290 72.840 ;
        RECT 8.890 71.740 9.290 72.840 ;
        RECT 10.890 71.740 11.290 72.840 ;
        RECT 12.890 71.740 13.290 72.840 ;
        RECT 14.890 71.740 15.290 72.840 ;
        RECT 16.890 71.740 17.290 72.840 ;
        RECT 18.890 71.740 19.290 72.840 ;
        RECT 20.890 71.740 21.290 72.840 ;
        RECT 22.890 71.740 23.290 72.840 ;
        RECT 24.890 71.740 25.290 72.840 ;
        RECT 26.890 71.740 27.290 72.840 ;
        RECT 28.890 71.740 29.290 72.840 ;
        RECT 30.890 71.740 31.290 72.840 ;
        RECT 32.890 71.740 33.290 72.840 ;
        RECT 34.890 71.740 35.290 72.840 ;
        RECT 36.890 71.740 37.290 72.840 ;
        RECT 38.890 71.740 39.290 72.840 ;
        RECT 40.890 71.740 41.290 72.840 ;
        RECT 42.890 71.740 43.290 72.840 ;
        RECT 44.890 71.740 45.290 72.840 ;
        RECT 46.890 71.740 47.290 72.840 ;
        RECT 48.890 71.740 49.290 72.840 ;
        RECT 50.890 71.740 51.290 72.840 ;
        RECT 52.890 71.740 53.290 72.840 ;
        RECT 54.890 71.740 55.290 72.840 ;
        RECT 56.890 71.740 57.290 72.840 ;
        RECT 58.890 71.740 59.290 72.840 ;
        RECT 60.890 71.740 61.290 72.840 ;
        RECT 62.890 71.740 63.290 72.840 ;
        RECT 64.890 71.740 65.290 72.840 ;
        RECT 66.890 71.740 67.290 72.840 ;
        RECT 68.890 71.740 69.290 72.840 ;
        RECT 70.890 71.740 71.290 72.840 ;
        RECT 72.890 71.740 73.290 72.840 ;
        RECT 6.890 69.890 7.290 70.990 ;
        RECT 8.890 69.890 9.290 70.990 ;
        RECT 10.890 69.890 11.290 70.990 ;
        RECT 12.890 69.890 13.290 70.990 ;
        RECT 14.890 69.890 15.290 70.990 ;
        RECT 16.890 69.890 17.290 70.990 ;
        RECT 18.890 69.890 19.290 70.990 ;
        RECT 20.890 69.890 21.290 70.990 ;
        RECT 22.890 69.890 23.290 70.990 ;
        RECT 24.890 69.890 25.290 70.990 ;
        RECT 26.890 69.890 27.290 70.990 ;
        RECT 28.890 69.890 29.290 70.990 ;
        RECT 30.890 69.890 31.290 70.990 ;
        RECT 32.890 69.890 33.290 70.990 ;
        RECT 34.890 69.890 35.290 70.990 ;
        RECT 36.890 69.890 37.290 70.990 ;
        RECT 38.890 69.890 39.290 70.990 ;
        RECT 40.890 69.890 41.290 70.990 ;
        RECT 42.890 69.890 43.290 70.990 ;
        RECT 44.890 69.890 45.290 70.990 ;
        RECT 46.890 69.890 47.290 70.990 ;
        RECT 48.890 69.890 49.290 70.990 ;
        RECT 50.890 69.890 51.290 70.990 ;
        RECT 52.890 69.890 53.290 70.990 ;
        RECT 54.890 69.890 55.290 70.990 ;
        RECT 56.890 69.890 57.290 70.990 ;
        RECT 58.890 69.890 59.290 70.990 ;
        RECT 60.890 69.890 61.290 70.990 ;
        RECT 62.890 69.890 63.290 70.990 ;
        RECT 64.890 69.890 65.290 70.990 ;
        RECT 66.890 69.890 67.290 70.990 ;
        RECT 68.890 69.890 69.290 70.990 ;
        RECT 70.890 69.890 71.290 70.990 ;
        RECT 72.890 69.890 73.290 70.990 ;
        RECT 6.890 68.040 7.290 69.140 ;
        RECT 8.890 68.040 9.290 69.140 ;
        RECT 10.890 68.040 11.290 69.140 ;
        RECT 12.890 68.040 13.290 69.140 ;
        RECT 14.890 68.040 15.290 69.140 ;
        RECT 16.890 68.040 17.290 69.140 ;
        RECT 18.890 68.040 19.290 69.140 ;
        RECT 20.890 68.040 21.290 69.140 ;
        RECT 22.890 68.040 23.290 69.140 ;
        RECT 24.890 68.040 25.290 69.140 ;
        RECT 26.890 68.040 27.290 69.140 ;
        RECT 28.890 68.040 29.290 69.140 ;
        RECT 30.890 68.040 31.290 69.140 ;
        RECT 32.890 68.040 33.290 69.140 ;
        RECT 34.890 68.040 35.290 69.140 ;
        RECT 36.890 68.040 37.290 69.140 ;
        RECT 38.890 68.040 39.290 69.140 ;
        RECT 40.890 68.040 41.290 69.140 ;
        RECT 42.890 68.040 43.290 69.140 ;
        RECT 44.890 68.040 45.290 69.140 ;
        RECT 46.890 68.040 47.290 69.140 ;
        RECT 48.890 68.040 49.290 69.140 ;
        RECT 50.890 68.040 51.290 69.140 ;
        RECT 52.890 68.040 53.290 69.140 ;
        RECT 54.890 68.040 55.290 69.140 ;
        RECT 56.890 68.040 57.290 69.140 ;
        RECT 58.890 68.040 59.290 69.140 ;
        RECT 60.890 68.040 61.290 69.140 ;
        RECT 62.890 68.040 63.290 69.140 ;
        RECT 64.890 68.040 65.290 69.140 ;
        RECT 66.890 68.040 67.290 69.140 ;
        RECT 68.890 68.040 69.290 69.140 ;
        RECT 70.890 68.040 71.290 69.140 ;
        RECT 72.890 68.040 73.290 69.140 ;
        RECT 6.890 66.190 7.290 67.290 ;
        RECT 8.890 66.190 9.290 67.290 ;
        RECT 10.890 66.190 11.290 67.290 ;
        RECT 12.890 66.190 13.290 67.290 ;
        RECT 14.890 66.190 15.290 67.290 ;
        RECT 16.890 66.190 17.290 67.290 ;
        RECT 18.890 66.190 19.290 67.290 ;
        RECT 20.890 66.190 21.290 67.290 ;
        RECT 22.890 66.190 23.290 67.290 ;
        RECT 24.890 66.190 25.290 67.290 ;
        RECT 26.890 66.190 27.290 67.290 ;
        RECT 28.890 66.190 29.290 67.290 ;
        RECT 30.890 66.190 31.290 67.290 ;
        RECT 32.890 66.190 33.290 67.290 ;
        RECT 34.890 66.190 35.290 67.290 ;
        RECT 36.890 66.190 37.290 67.290 ;
        RECT 38.890 66.190 39.290 67.290 ;
        RECT 40.890 66.190 41.290 67.290 ;
        RECT 42.890 66.190 43.290 67.290 ;
        RECT 44.890 66.190 45.290 67.290 ;
        RECT 46.890 66.190 47.290 67.290 ;
        RECT 48.890 66.190 49.290 67.290 ;
        RECT 50.890 66.190 51.290 67.290 ;
        RECT 52.890 66.190 53.290 67.290 ;
        RECT 54.890 66.190 55.290 67.290 ;
        RECT 56.890 66.190 57.290 67.290 ;
        RECT 58.890 66.190 59.290 67.290 ;
        RECT 60.890 66.190 61.290 67.290 ;
        RECT 62.890 66.190 63.290 67.290 ;
        RECT 64.890 66.190 65.290 67.290 ;
        RECT 66.890 66.190 67.290 67.290 ;
        RECT 68.890 66.190 69.290 67.290 ;
        RECT 70.890 66.190 71.290 67.290 ;
        RECT 72.890 66.190 73.290 67.290 ;
        RECT 6.890 64.340 7.290 65.440 ;
        RECT 8.890 64.340 9.290 65.440 ;
        RECT 10.890 64.340 11.290 65.440 ;
        RECT 12.890 64.340 13.290 65.440 ;
        RECT 14.890 64.340 15.290 65.440 ;
        RECT 16.890 64.340 17.290 65.440 ;
        RECT 18.890 64.340 19.290 65.440 ;
        RECT 20.890 64.340 21.290 65.440 ;
        RECT 22.890 64.340 23.290 65.440 ;
        RECT 24.890 64.340 25.290 65.440 ;
        RECT 26.890 64.340 27.290 65.440 ;
        RECT 28.890 64.340 29.290 65.440 ;
        RECT 30.890 64.340 31.290 65.440 ;
        RECT 32.890 64.340 33.290 65.440 ;
        RECT 34.890 64.340 35.290 65.440 ;
        RECT 36.890 64.340 37.290 65.440 ;
        RECT 38.890 64.340 39.290 65.440 ;
        RECT 40.890 64.340 41.290 65.440 ;
        RECT 42.890 64.340 43.290 65.440 ;
        RECT 44.890 64.340 45.290 65.440 ;
        RECT 46.890 64.340 47.290 65.440 ;
        RECT 48.890 64.340 49.290 65.440 ;
        RECT 50.890 64.340 51.290 65.440 ;
        RECT 52.890 64.340 53.290 65.440 ;
        RECT 54.890 64.340 55.290 65.440 ;
        RECT 56.890 64.340 57.290 65.440 ;
        RECT 58.890 64.340 59.290 65.440 ;
        RECT 60.890 64.340 61.290 65.440 ;
        RECT 62.890 64.340 63.290 65.440 ;
        RECT 64.890 64.340 65.290 65.440 ;
        RECT 66.890 64.340 67.290 65.440 ;
        RECT 68.890 64.340 69.290 65.440 ;
        RECT 70.890 64.340 71.290 65.440 ;
        RECT 72.890 64.340 73.290 65.440 ;
        RECT 6.890 62.490 7.290 63.590 ;
        RECT 8.890 62.490 9.290 63.590 ;
        RECT 10.890 62.490 11.290 63.590 ;
        RECT 12.890 62.490 13.290 63.590 ;
        RECT 14.890 62.490 15.290 63.590 ;
        RECT 16.890 62.490 17.290 63.590 ;
        RECT 18.890 62.490 19.290 63.590 ;
        RECT 20.890 62.490 21.290 63.590 ;
        RECT 22.890 62.490 23.290 63.590 ;
        RECT 24.890 62.490 25.290 63.590 ;
        RECT 26.890 62.490 27.290 63.590 ;
        RECT 28.890 62.490 29.290 63.590 ;
        RECT 30.890 62.490 31.290 63.590 ;
        RECT 32.890 62.490 33.290 63.590 ;
        RECT 34.890 62.490 35.290 63.590 ;
        RECT 36.890 62.490 37.290 63.590 ;
        RECT 38.890 62.490 39.290 63.590 ;
        RECT 40.890 62.490 41.290 63.590 ;
        RECT 42.890 62.490 43.290 63.590 ;
        RECT 44.890 62.490 45.290 63.590 ;
        RECT 46.890 62.490 47.290 63.590 ;
        RECT 48.890 62.490 49.290 63.590 ;
        RECT 50.890 62.490 51.290 63.590 ;
        RECT 52.890 62.490 53.290 63.590 ;
        RECT 54.890 62.490 55.290 63.590 ;
        RECT 56.890 62.490 57.290 63.590 ;
        RECT 58.890 62.490 59.290 63.590 ;
        RECT 60.890 62.490 61.290 63.590 ;
        RECT 62.890 62.490 63.290 63.590 ;
        RECT 64.890 62.490 65.290 63.590 ;
        RECT 66.890 62.490 67.290 63.590 ;
        RECT 68.890 62.490 69.290 63.590 ;
        RECT 70.890 62.490 71.290 63.590 ;
        RECT 72.890 62.490 73.290 63.590 ;
        RECT 6.890 60.640 7.290 61.740 ;
        RECT 8.890 60.640 9.290 61.740 ;
        RECT 10.890 60.640 11.290 61.740 ;
        RECT 12.890 60.640 13.290 61.740 ;
        RECT 14.890 60.640 15.290 61.740 ;
        RECT 16.890 60.640 17.290 61.740 ;
        RECT 18.890 60.640 19.290 61.740 ;
        RECT 20.890 60.640 21.290 61.740 ;
        RECT 22.890 60.640 23.290 61.740 ;
        RECT 24.890 60.640 25.290 61.740 ;
        RECT 26.890 60.640 27.290 61.740 ;
        RECT 28.890 60.640 29.290 61.740 ;
        RECT 30.890 60.640 31.290 61.740 ;
        RECT 32.890 60.640 33.290 61.740 ;
        RECT 34.890 60.640 35.290 61.740 ;
        RECT 36.890 60.640 37.290 61.740 ;
        RECT 38.890 60.640 39.290 61.740 ;
        RECT 40.890 60.640 41.290 61.740 ;
        RECT 42.890 60.640 43.290 61.740 ;
        RECT 44.890 60.640 45.290 61.740 ;
        RECT 46.890 60.640 47.290 61.740 ;
        RECT 48.890 60.640 49.290 61.740 ;
        RECT 50.890 60.640 51.290 61.740 ;
        RECT 52.890 60.640 53.290 61.740 ;
        RECT 54.890 60.640 55.290 61.740 ;
        RECT 56.890 60.640 57.290 61.740 ;
        RECT 58.890 60.640 59.290 61.740 ;
        RECT 60.890 60.640 61.290 61.740 ;
        RECT 62.890 60.640 63.290 61.740 ;
        RECT 64.890 60.640 65.290 61.740 ;
        RECT 66.890 60.640 67.290 61.740 ;
        RECT 68.890 60.640 69.290 61.740 ;
        RECT 70.890 60.640 71.290 61.740 ;
        RECT 72.890 60.640 73.290 61.740 ;
        RECT 6.890 58.790 7.290 59.890 ;
        RECT 8.890 58.790 9.290 59.890 ;
        RECT 10.890 58.790 11.290 59.890 ;
        RECT 12.890 58.790 13.290 59.890 ;
        RECT 14.890 58.790 15.290 59.890 ;
        RECT 16.890 58.790 17.290 59.890 ;
        RECT 18.890 58.790 19.290 59.890 ;
        RECT 20.890 58.790 21.290 59.890 ;
        RECT 22.890 58.790 23.290 59.890 ;
        RECT 24.890 58.790 25.290 59.890 ;
        RECT 26.890 58.790 27.290 59.890 ;
        RECT 28.890 58.790 29.290 59.890 ;
        RECT 30.890 58.790 31.290 59.890 ;
        RECT 32.890 58.790 33.290 59.890 ;
        RECT 34.890 58.790 35.290 59.890 ;
        RECT 36.890 58.790 37.290 59.890 ;
        RECT 38.890 58.790 39.290 59.890 ;
        RECT 40.890 58.790 41.290 59.890 ;
        RECT 42.890 58.790 43.290 59.890 ;
        RECT 44.890 58.790 45.290 59.890 ;
        RECT 46.890 58.790 47.290 59.890 ;
        RECT 48.890 58.790 49.290 59.890 ;
        RECT 50.890 58.790 51.290 59.890 ;
        RECT 52.890 58.790 53.290 59.890 ;
        RECT 54.890 58.790 55.290 59.890 ;
        RECT 56.890 58.790 57.290 59.890 ;
        RECT 58.890 58.790 59.290 59.890 ;
        RECT 60.890 58.790 61.290 59.890 ;
        RECT 62.890 58.790 63.290 59.890 ;
        RECT 64.890 58.790 65.290 59.890 ;
        RECT 66.890 58.790 67.290 59.890 ;
        RECT 68.890 58.790 69.290 59.890 ;
        RECT 70.890 58.790 71.290 59.890 ;
        RECT 72.890 58.790 73.290 59.890 ;
        RECT 6.890 56.940 7.290 58.040 ;
        RECT 8.890 56.940 9.290 58.040 ;
        RECT 10.890 56.940 11.290 58.040 ;
        RECT 12.890 56.940 13.290 58.040 ;
        RECT 14.890 56.940 15.290 58.040 ;
        RECT 16.890 56.940 17.290 58.040 ;
        RECT 18.890 56.940 19.290 58.040 ;
        RECT 20.890 56.940 21.290 58.040 ;
        RECT 22.890 56.940 23.290 58.040 ;
        RECT 24.890 56.940 25.290 58.040 ;
        RECT 26.890 56.940 27.290 58.040 ;
        RECT 28.890 56.940 29.290 58.040 ;
        RECT 30.890 56.940 31.290 58.040 ;
        RECT 32.890 56.940 33.290 58.040 ;
        RECT 34.890 56.940 35.290 58.040 ;
        RECT 36.890 56.940 37.290 58.040 ;
        RECT 38.890 56.940 39.290 58.040 ;
        RECT 40.890 56.940 41.290 58.040 ;
        RECT 42.890 56.940 43.290 58.040 ;
        RECT 44.890 56.940 45.290 58.040 ;
        RECT 46.890 56.940 47.290 58.040 ;
        RECT 48.890 56.940 49.290 58.040 ;
        RECT 50.890 56.940 51.290 58.040 ;
        RECT 52.890 56.940 53.290 58.040 ;
        RECT 54.890 56.940 55.290 58.040 ;
        RECT 56.890 56.940 57.290 58.040 ;
        RECT 58.890 56.940 59.290 58.040 ;
        RECT 60.890 56.940 61.290 58.040 ;
        RECT 62.890 56.940 63.290 58.040 ;
        RECT 64.890 56.940 65.290 58.040 ;
        RECT 66.890 56.940 67.290 58.040 ;
        RECT 68.890 56.940 69.290 58.040 ;
        RECT 70.890 56.940 71.290 58.040 ;
        RECT 72.890 56.940 73.290 58.040 ;
        RECT 6.890 55.090 7.290 56.190 ;
        RECT 8.890 55.090 9.290 56.190 ;
        RECT 10.890 55.090 11.290 56.190 ;
        RECT 12.890 55.090 13.290 56.190 ;
        RECT 14.890 55.090 15.290 56.190 ;
        RECT 16.890 55.090 17.290 56.190 ;
        RECT 18.890 55.090 19.290 56.190 ;
        RECT 20.890 55.090 21.290 56.190 ;
        RECT 22.890 55.090 23.290 56.190 ;
        RECT 24.890 55.090 25.290 56.190 ;
        RECT 26.890 55.090 27.290 56.190 ;
        RECT 28.890 55.090 29.290 56.190 ;
        RECT 30.890 55.090 31.290 56.190 ;
        RECT 32.890 55.090 33.290 56.190 ;
        RECT 34.890 55.090 35.290 56.190 ;
        RECT 36.890 55.090 37.290 56.190 ;
        RECT 38.890 55.090 39.290 56.190 ;
        RECT 40.890 55.090 41.290 56.190 ;
        RECT 42.890 55.090 43.290 56.190 ;
        RECT 44.890 55.090 45.290 56.190 ;
        RECT 46.890 55.090 47.290 56.190 ;
        RECT 48.890 55.090 49.290 56.190 ;
        RECT 50.890 55.090 51.290 56.190 ;
        RECT 52.890 55.090 53.290 56.190 ;
        RECT 54.890 55.090 55.290 56.190 ;
        RECT 56.890 55.090 57.290 56.190 ;
        RECT 58.890 55.090 59.290 56.190 ;
        RECT 60.890 55.090 61.290 56.190 ;
        RECT 62.890 55.090 63.290 56.190 ;
        RECT 64.890 55.090 65.290 56.190 ;
        RECT 66.890 55.090 67.290 56.190 ;
        RECT 68.890 55.090 69.290 56.190 ;
        RECT 70.890 55.090 71.290 56.190 ;
        RECT 72.890 55.090 73.290 56.190 ;
        RECT 6.890 53.240 7.290 54.340 ;
        RECT 8.890 53.240 9.290 54.340 ;
        RECT 10.890 53.240 11.290 54.340 ;
        RECT 12.890 53.240 13.290 54.340 ;
        RECT 14.890 53.240 15.290 54.340 ;
        RECT 16.890 53.240 17.290 54.340 ;
        RECT 18.890 53.240 19.290 54.340 ;
        RECT 20.890 53.240 21.290 54.340 ;
        RECT 22.890 53.240 23.290 54.340 ;
        RECT 24.890 53.240 25.290 54.340 ;
        RECT 26.890 53.240 27.290 54.340 ;
        RECT 28.890 53.240 29.290 54.340 ;
        RECT 30.890 53.240 31.290 54.340 ;
        RECT 32.890 53.240 33.290 54.340 ;
        RECT 34.890 53.240 35.290 54.340 ;
        RECT 36.890 53.240 37.290 54.340 ;
        RECT 38.890 53.240 39.290 54.340 ;
        RECT 40.890 53.240 41.290 54.340 ;
        RECT 42.890 53.240 43.290 54.340 ;
        RECT 44.890 53.240 45.290 54.340 ;
        RECT 46.890 53.240 47.290 54.340 ;
        RECT 48.890 53.240 49.290 54.340 ;
        RECT 50.890 53.240 51.290 54.340 ;
        RECT 52.890 53.240 53.290 54.340 ;
        RECT 54.890 53.240 55.290 54.340 ;
        RECT 56.890 53.240 57.290 54.340 ;
        RECT 58.890 53.240 59.290 54.340 ;
        RECT 60.890 53.240 61.290 54.340 ;
        RECT 62.890 53.240 63.290 54.340 ;
        RECT 64.890 53.240 65.290 54.340 ;
        RECT 66.890 53.240 67.290 54.340 ;
        RECT 68.890 53.240 69.290 54.340 ;
        RECT 70.890 53.240 71.290 54.340 ;
        RECT 72.890 53.240 73.290 54.340 ;
        RECT 6.890 51.390 7.290 52.490 ;
        RECT 8.890 51.390 9.290 52.490 ;
        RECT 10.890 51.390 11.290 52.490 ;
        RECT 12.890 51.390 13.290 52.490 ;
        RECT 14.890 51.390 15.290 52.490 ;
        RECT 16.890 51.390 17.290 52.490 ;
        RECT 18.890 51.390 19.290 52.490 ;
        RECT 20.890 51.390 21.290 52.490 ;
        RECT 22.890 51.390 23.290 52.490 ;
        RECT 24.890 51.390 25.290 52.490 ;
        RECT 26.890 51.390 27.290 52.490 ;
        RECT 28.890 51.390 29.290 52.490 ;
        RECT 30.890 51.390 31.290 52.490 ;
        RECT 32.890 51.390 33.290 52.490 ;
        RECT 34.890 51.390 35.290 52.490 ;
        RECT 36.890 51.390 37.290 52.490 ;
        RECT 38.890 51.390 39.290 52.490 ;
        RECT 40.890 51.390 41.290 52.490 ;
        RECT 42.890 51.390 43.290 52.490 ;
        RECT 44.890 51.390 45.290 52.490 ;
        RECT 46.890 51.390 47.290 52.490 ;
        RECT 48.890 51.390 49.290 52.490 ;
        RECT 50.890 51.390 51.290 52.490 ;
        RECT 52.890 51.390 53.290 52.490 ;
        RECT 54.890 51.390 55.290 52.490 ;
        RECT 56.890 51.390 57.290 52.490 ;
        RECT 58.890 51.390 59.290 52.490 ;
        RECT 60.890 51.390 61.290 52.490 ;
        RECT 62.890 51.390 63.290 52.490 ;
        RECT 64.890 51.390 65.290 52.490 ;
        RECT 66.890 51.390 67.290 52.490 ;
        RECT 68.890 51.390 69.290 52.490 ;
        RECT 70.890 51.390 71.290 52.490 ;
        RECT 72.890 51.390 73.290 52.490 ;
        RECT 6.890 49.540 7.290 50.640 ;
        RECT 8.890 49.540 9.290 50.640 ;
        RECT 10.890 49.540 11.290 50.640 ;
        RECT 12.890 49.540 13.290 50.640 ;
        RECT 14.890 49.540 15.290 50.640 ;
        RECT 16.890 49.540 17.290 50.640 ;
        RECT 18.890 49.540 19.290 50.640 ;
        RECT 20.890 49.540 21.290 50.640 ;
        RECT 22.890 49.540 23.290 50.640 ;
        RECT 24.890 49.540 25.290 50.640 ;
        RECT 26.890 49.540 27.290 50.640 ;
        RECT 28.890 49.540 29.290 50.640 ;
        RECT 30.890 49.540 31.290 50.640 ;
        RECT 32.890 49.540 33.290 50.640 ;
        RECT 34.890 49.540 35.290 50.640 ;
        RECT 36.890 49.540 37.290 50.640 ;
        RECT 38.890 49.540 39.290 50.640 ;
        RECT 40.890 49.540 41.290 50.640 ;
        RECT 42.890 49.540 43.290 50.640 ;
        RECT 44.890 49.540 45.290 50.640 ;
        RECT 46.890 49.540 47.290 50.640 ;
        RECT 48.890 49.540 49.290 50.640 ;
        RECT 50.890 49.540 51.290 50.640 ;
        RECT 52.890 49.540 53.290 50.640 ;
        RECT 54.890 49.540 55.290 50.640 ;
        RECT 56.890 49.540 57.290 50.640 ;
        RECT 58.890 49.540 59.290 50.640 ;
        RECT 60.890 49.540 61.290 50.640 ;
        RECT 62.890 49.540 63.290 50.640 ;
        RECT 64.890 49.540 65.290 50.640 ;
        RECT 66.890 49.540 67.290 50.640 ;
        RECT 68.890 49.540 69.290 50.640 ;
        RECT 70.890 49.540 71.290 50.640 ;
        RECT 72.890 49.540 73.290 50.640 ;
        RECT 6.890 47.690 7.290 48.790 ;
        RECT 8.890 47.690 9.290 48.790 ;
        RECT 10.890 47.690 11.290 48.790 ;
        RECT 12.890 47.690 13.290 48.790 ;
        RECT 14.890 47.690 15.290 48.790 ;
        RECT 16.890 47.690 17.290 48.790 ;
        RECT 18.890 47.690 19.290 48.790 ;
        RECT 20.890 47.690 21.290 48.790 ;
        RECT 22.890 47.690 23.290 48.790 ;
        RECT 24.890 47.690 25.290 48.790 ;
        RECT 26.890 47.690 27.290 48.790 ;
        RECT 28.890 47.690 29.290 48.790 ;
        RECT 30.890 47.690 31.290 48.790 ;
        RECT 32.890 47.690 33.290 48.790 ;
        RECT 34.890 47.690 35.290 48.790 ;
        RECT 36.890 47.690 37.290 48.790 ;
        RECT 38.890 47.690 39.290 48.790 ;
        RECT 40.890 47.690 41.290 48.790 ;
        RECT 42.890 47.690 43.290 48.790 ;
        RECT 44.890 47.690 45.290 48.790 ;
        RECT 46.890 47.690 47.290 48.790 ;
        RECT 48.890 47.690 49.290 48.790 ;
        RECT 50.890 47.690 51.290 48.790 ;
        RECT 52.890 47.690 53.290 48.790 ;
        RECT 54.890 47.690 55.290 48.790 ;
        RECT 56.890 47.690 57.290 48.790 ;
        RECT 58.890 47.690 59.290 48.790 ;
        RECT 60.890 47.690 61.290 48.790 ;
        RECT 62.890 47.690 63.290 48.790 ;
        RECT 64.890 47.690 65.290 48.790 ;
        RECT 66.890 47.690 67.290 48.790 ;
        RECT 68.890 47.690 69.290 48.790 ;
        RECT 70.890 47.690 71.290 48.790 ;
        RECT 72.890 47.690 73.290 48.790 ;
        RECT 6.890 45.840 7.290 46.940 ;
        RECT 8.890 45.840 9.290 46.940 ;
        RECT 10.890 45.840 11.290 46.940 ;
        RECT 12.890 45.840 13.290 46.940 ;
        RECT 14.890 45.840 15.290 46.940 ;
        RECT 16.890 45.840 17.290 46.940 ;
        RECT 18.890 45.840 19.290 46.940 ;
        RECT 20.890 45.840 21.290 46.940 ;
        RECT 22.890 45.840 23.290 46.940 ;
        RECT 24.890 45.840 25.290 46.940 ;
        RECT 26.890 45.840 27.290 46.940 ;
        RECT 28.890 45.840 29.290 46.940 ;
        RECT 30.890 45.840 31.290 46.940 ;
        RECT 32.890 45.840 33.290 46.940 ;
        RECT 34.890 45.840 35.290 46.940 ;
        RECT 36.890 45.840 37.290 46.940 ;
        RECT 38.890 45.840 39.290 46.940 ;
        RECT 40.890 45.840 41.290 46.940 ;
        RECT 42.890 45.840 43.290 46.940 ;
        RECT 44.890 45.840 45.290 46.940 ;
        RECT 46.890 45.840 47.290 46.940 ;
        RECT 48.890 45.840 49.290 46.940 ;
        RECT 50.890 45.840 51.290 46.940 ;
        RECT 52.890 45.840 53.290 46.940 ;
        RECT 54.890 45.840 55.290 46.940 ;
        RECT 56.890 45.840 57.290 46.940 ;
        RECT 58.890 45.840 59.290 46.940 ;
        RECT 60.890 45.840 61.290 46.940 ;
        RECT 62.890 45.840 63.290 46.940 ;
        RECT 64.890 45.840 65.290 46.940 ;
        RECT 66.890 45.840 67.290 46.940 ;
        RECT 68.890 45.840 69.290 46.940 ;
        RECT 70.890 45.840 71.290 46.940 ;
        RECT 72.890 45.840 73.290 46.940 ;
        RECT 6.890 43.990 7.290 45.090 ;
        RECT 8.890 43.990 9.290 45.090 ;
        RECT 10.890 43.990 11.290 45.090 ;
        RECT 12.890 43.990 13.290 45.090 ;
        RECT 14.890 43.990 15.290 45.090 ;
        RECT 16.890 43.990 17.290 45.090 ;
        RECT 18.890 43.990 19.290 45.090 ;
        RECT 20.890 43.990 21.290 45.090 ;
        RECT 22.890 43.990 23.290 45.090 ;
        RECT 24.890 43.990 25.290 45.090 ;
        RECT 26.890 43.990 27.290 45.090 ;
        RECT 28.890 43.990 29.290 45.090 ;
        RECT 30.890 43.990 31.290 45.090 ;
        RECT 32.890 43.990 33.290 45.090 ;
        RECT 34.890 43.990 35.290 45.090 ;
        RECT 36.890 43.990 37.290 45.090 ;
        RECT 38.890 43.990 39.290 45.090 ;
        RECT 40.890 43.990 41.290 45.090 ;
        RECT 42.890 43.990 43.290 45.090 ;
        RECT 44.890 43.990 45.290 45.090 ;
        RECT 46.890 43.990 47.290 45.090 ;
        RECT 48.890 43.990 49.290 45.090 ;
        RECT 50.890 43.990 51.290 45.090 ;
        RECT 52.890 43.990 53.290 45.090 ;
        RECT 54.890 43.990 55.290 45.090 ;
        RECT 56.890 43.990 57.290 45.090 ;
        RECT 58.890 43.990 59.290 45.090 ;
        RECT 60.890 43.990 61.290 45.090 ;
        RECT 62.890 43.990 63.290 45.090 ;
        RECT 64.890 43.990 65.290 45.090 ;
        RECT 66.890 43.990 67.290 45.090 ;
        RECT 68.890 43.990 69.290 45.090 ;
        RECT 70.890 43.990 71.290 45.090 ;
        RECT 72.890 43.990 73.290 45.090 ;
        RECT 6.890 42.140 7.290 43.240 ;
        RECT 8.890 42.140 9.290 43.240 ;
        RECT 10.890 42.140 11.290 43.240 ;
        RECT 12.890 42.140 13.290 43.240 ;
        RECT 14.890 42.140 15.290 43.240 ;
        RECT 16.890 42.140 17.290 43.240 ;
        RECT 18.890 42.140 19.290 43.240 ;
        RECT 20.890 42.140 21.290 43.240 ;
        RECT 22.890 42.140 23.290 43.240 ;
        RECT 24.890 42.140 25.290 43.240 ;
        RECT 26.890 42.140 27.290 43.240 ;
        RECT 28.890 42.140 29.290 43.240 ;
        RECT 30.890 42.140 31.290 43.240 ;
        RECT 32.890 42.140 33.290 43.240 ;
        RECT 34.890 42.140 35.290 43.240 ;
        RECT 36.890 42.140 37.290 43.240 ;
        RECT 38.890 42.140 39.290 43.240 ;
        RECT 40.890 42.140 41.290 43.240 ;
        RECT 42.890 42.140 43.290 43.240 ;
        RECT 44.890 42.140 45.290 43.240 ;
        RECT 46.890 42.140 47.290 43.240 ;
        RECT 48.890 42.140 49.290 43.240 ;
        RECT 50.890 42.140 51.290 43.240 ;
        RECT 52.890 42.140 53.290 43.240 ;
        RECT 54.890 42.140 55.290 43.240 ;
        RECT 56.890 42.140 57.290 43.240 ;
        RECT 58.890 42.140 59.290 43.240 ;
        RECT 60.890 42.140 61.290 43.240 ;
        RECT 62.890 42.140 63.290 43.240 ;
        RECT 64.890 42.140 65.290 43.240 ;
        RECT 66.890 42.140 67.290 43.240 ;
        RECT 68.890 42.140 69.290 43.240 ;
        RECT 70.890 42.140 71.290 43.240 ;
        RECT 72.890 42.140 73.290 43.240 ;
        RECT 6.890 40.290 7.290 41.390 ;
        RECT 8.890 40.290 9.290 41.390 ;
        RECT 10.890 40.290 11.290 41.390 ;
        RECT 12.890 40.290 13.290 41.390 ;
        RECT 14.890 40.290 15.290 41.390 ;
        RECT 16.890 40.290 17.290 41.390 ;
        RECT 18.890 40.290 19.290 41.390 ;
        RECT 20.890 40.290 21.290 41.390 ;
        RECT 22.890 40.290 23.290 41.390 ;
        RECT 24.890 40.290 25.290 41.390 ;
        RECT 26.890 40.290 27.290 41.390 ;
        RECT 28.890 40.290 29.290 41.390 ;
        RECT 30.890 40.290 31.290 41.390 ;
        RECT 32.890 40.290 33.290 41.390 ;
        RECT 34.890 40.290 35.290 41.390 ;
        RECT 36.890 40.290 37.290 41.390 ;
        RECT 38.890 40.290 39.290 41.390 ;
        RECT 40.890 40.290 41.290 41.390 ;
        RECT 42.890 40.290 43.290 41.390 ;
        RECT 44.890 40.290 45.290 41.390 ;
        RECT 46.890 40.290 47.290 41.390 ;
        RECT 48.890 40.290 49.290 41.390 ;
        RECT 50.890 40.290 51.290 41.390 ;
        RECT 52.890 40.290 53.290 41.390 ;
        RECT 54.890 40.290 55.290 41.390 ;
        RECT 56.890 40.290 57.290 41.390 ;
        RECT 58.890 40.290 59.290 41.390 ;
        RECT 60.890 40.290 61.290 41.390 ;
        RECT 62.890 40.290 63.290 41.390 ;
        RECT 64.890 40.290 65.290 41.390 ;
        RECT 66.890 40.290 67.290 41.390 ;
        RECT 68.890 40.290 69.290 41.390 ;
        RECT 70.890 40.290 71.290 41.390 ;
        RECT 72.890 40.290 73.290 41.390 ;
        RECT 6.890 38.440 7.290 39.540 ;
        RECT 8.890 38.440 9.290 39.540 ;
        RECT 10.890 38.440 11.290 39.540 ;
        RECT 12.890 38.440 13.290 39.540 ;
        RECT 14.890 38.440 15.290 39.540 ;
        RECT 16.890 38.440 17.290 39.540 ;
        RECT 18.890 38.440 19.290 39.540 ;
        RECT 20.890 38.440 21.290 39.540 ;
        RECT 22.890 38.440 23.290 39.540 ;
        RECT 24.890 38.440 25.290 39.540 ;
        RECT 26.890 38.440 27.290 39.540 ;
        RECT 28.890 38.440 29.290 39.540 ;
        RECT 30.890 38.440 31.290 39.540 ;
        RECT 32.890 38.440 33.290 39.540 ;
        RECT 34.890 38.440 35.290 39.540 ;
        RECT 36.890 38.440 37.290 39.540 ;
        RECT 38.890 38.440 39.290 39.540 ;
        RECT 40.890 38.440 41.290 39.540 ;
        RECT 42.890 38.440 43.290 39.540 ;
        RECT 44.890 38.440 45.290 39.540 ;
        RECT 46.890 38.440 47.290 39.540 ;
        RECT 48.890 38.440 49.290 39.540 ;
        RECT 50.890 38.440 51.290 39.540 ;
        RECT 52.890 38.440 53.290 39.540 ;
        RECT 54.890 38.440 55.290 39.540 ;
        RECT 56.890 38.440 57.290 39.540 ;
        RECT 58.890 38.440 59.290 39.540 ;
        RECT 60.890 38.440 61.290 39.540 ;
        RECT 62.890 38.440 63.290 39.540 ;
        RECT 64.890 38.440 65.290 39.540 ;
        RECT 66.890 38.440 67.290 39.540 ;
        RECT 68.890 38.440 69.290 39.540 ;
        RECT 70.890 38.440 71.290 39.540 ;
        RECT 72.890 38.440 73.290 39.540 ;
        RECT 6.890 36.590 7.290 37.690 ;
        RECT 8.890 36.590 9.290 37.690 ;
        RECT 10.890 36.590 11.290 37.690 ;
        RECT 12.890 36.590 13.290 37.690 ;
        RECT 14.890 36.590 15.290 37.690 ;
        RECT 16.890 36.590 17.290 37.690 ;
        RECT 18.890 36.590 19.290 37.690 ;
        RECT 20.890 36.590 21.290 37.690 ;
        RECT 22.890 36.590 23.290 37.690 ;
        RECT 24.890 36.590 25.290 37.690 ;
        RECT 26.890 36.590 27.290 37.690 ;
        RECT 28.890 36.590 29.290 37.690 ;
        RECT 30.890 36.590 31.290 37.690 ;
        RECT 32.890 36.590 33.290 37.690 ;
        RECT 34.890 36.590 35.290 37.690 ;
        RECT 36.890 36.590 37.290 37.690 ;
        RECT 38.890 36.590 39.290 37.690 ;
        RECT 40.890 36.590 41.290 37.690 ;
        RECT 42.890 36.590 43.290 37.690 ;
        RECT 44.890 36.590 45.290 37.690 ;
        RECT 46.890 36.590 47.290 37.690 ;
        RECT 48.890 36.590 49.290 37.690 ;
        RECT 50.890 36.590 51.290 37.690 ;
        RECT 52.890 36.590 53.290 37.690 ;
        RECT 54.890 36.590 55.290 37.690 ;
        RECT 56.890 36.590 57.290 37.690 ;
        RECT 58.890 36.590 59.290 37.690 ;
        RECT 60.890 36.590 61.290 37.690 ;
        RECT 62.890 36.590 63.290 37.690 ;
        RECT 64.890 36.590 65.290 37.690 ;
        RECT 66.890 36.590 67.290 37.690 ;
        RECT 68.890 36.590 69.290 37.690 ;
        RECT 70.890 36.590 71.290 37.690 ;
        RECT 72.890 36.590 73.290 37.690 ;
        RECT 6.890 34.740 7.290 35.840 ;
        RECT 8.890 34.740 9.290 35.840 ;
        RECT 10.890 34.740 11.290 35.840 ;
        RECT 12.890 34.740 13.290 35.840 ;
        RECT 14.890 34.740 15.290 35.840 ;
        RECT 16.890 34.740 17.290 35.840 ;
        RECT 18.890 34.740 19.290 35.840 ;
        RECT 20.890 34.740 21.290 35.840 ;
        RECT 22.890 34.740 23.290 35.840 ;
        RECT 24.890 34.740 25.290 35.840 ;
        RECT 26.890 34.740 27.290 35.840 ;
        RECT 28.890 34.740 29.290 35.840 ;
        RECT 30.890 34.740 31.290 35.840 ;
        RECT 32.890 34.740 33.290 35.840 ;
        RECT 34.890 34.740 35.290 35.840 ;
        RECT 36.890 34.740 37.290 35.840 ;
        RECT 38.890 34.740 39.290 35.840 ;
        RECT 40.890 34.740 41.290 35.840 ;
        RECT 42.890 34.740 43.290 35.840 ;
        RECT 44.890 34.740 45.290 35.840 ;
        RECT 46.890 34.740 47.290 35.840 ;
        RECT 48.890 34.740 49.290 35.840 ;
        RECT 50.890 34.740 51.290 35.840 ;
        RECT 52.890 34.740 53.290 35.840 ;
        RECT 54.890 34.740 55.290 35.840 ;
        RECT 56.890 34.740 57.290 35.840 ;
        RECT 58.890 34.740 59.290 35.840 ;
        RECT 60.890 34.740 61.290 35.840 ;
        RECT 62.890 34.740 63.290 35.840 ;
        RECT 64.890 34.740 65.290 35.840 ;
        RECT 66.890 34.740 67.290 35.840 ;
        RECT 68.890 34.740 69.290 35.840 ;
        RECT 70.890 34.740 71.290 35.840 ;
        RECT 72.890 34.740 73.290 35.840 ;
        RECT 6.890 32.890 7.290 33.990 ;
        RECT 8.890 32.890 9.290 33.990 ;
        RECT 10.890 32.890 11.290 33.990 ;
        RECT 12.890 32.890 13.290 33.990 ;
        RECT 14.890 32.890 15.290 33.990 ;
        RECT 16.890 32.890 17.290 33.990 ;
        RECT 18.890 32.890 19.290 33.990 ;
        RECT 20.890 32.890 21.290 33.990 ;
        RECT 22.890 32.890 23.290 33.990 ;
        RECT 24.890 32.890 25.290 33.990 ;
        RECT 26.890 32.890 27.290 33.990 ;
        RECT 28.890 32.890 29.290 33.990 ;
        RECT 30.890 32.890 31.290 33.990 ;
        RECT 32.890 32.890 33.290 33.990 ;
        RECT 34.890 32.890 35.290 33.990 ;
        RECT 36.890 32.890 37.290 33.990 ;
        RECT 38.890 32.890 39.290 33.990 ;
        RECT 40.890 32.890 41.290 33.990 ;
        RECT 42.890 32.890 43.290 33.990 ;
        RECT 44.890 32.890 45.290 33.990 ;
        RECT 46.890 32.890 47.290 33.990 ;
        RECT 48.890 32.890 49.290 33.990 ;
        RECT 50.890 32.890 51.290 33.990 ;
        RECT 52.890 32.890 53.290 33.990 ;
        RECT 54.890 32.890 55.290 33.990 ;
        RECT 56.890 32.890 57.290 33.990 ;
        RECT 58.890 32.890 59.290 33.990 ;
        RECT 60.890 32.890 61.290 33.990 ;
        RECT 62.890 32.890 63.290 33.990 ;
        RECT 64.890 32.890 65.290 33.990 ;
        RECT 66.890 32.890 67.290 33.990 ;
        RECT 68.890 32.890 69.290 33.990 ;
        RECT 70.890 32.890 71.290 33.990 ;
        RECT 72.890 32.890 73.290 33.990 ;
        RECT 6.890 31.040 7.290 32.140 ;
        RECT 8.890 31.040 9.290 32.140 ;
        RECT 10.890 31.040 11.290 32.140 ;
        RECT 12.890 31.040 13.290 32.140 ;
        RECT 14.890 31.040 15.290 32.140 ;
        RECT 16.890 31.040 17.290 32.140 ;
        RECT 18.890 31.040 19.290 32.140 ;
        RECT 20.890 31.040 21.290 32.140 ;
        RECT 22.890 31.040 23.290 32.140 ;
        RECT 24.890 31.040 25.290 32.140 ;
        RECT 26.890 31.040 27.290 32.140 ;
        RECT 28.890 31.040 29.290 32.140 ;
        RECT 30.890 31.040 31.290 32.140 ;
        RECT 32.890 31.040 33.290 32.140 ;
        RECT 34.890 31.040 35.290 32.140 ;
        RECT 36.890 31.040 37.290 32.140 ;
        RECT 38.890 31.040 39.290 32.140 ;
        RECT 40.890 31.040 41.290 32.140 ;
        RECT 42.890 31.040 43.290 32.140 ;
        RECT 44.890 31.040 45.290 32.140 ;
        RECT 46.890 31.040 47.290 32.140 ;
        RECT 48.890 31.040 49.290 32.140 ;
        RECT 50.890 31.040 51.290 32.140 ;
        RECT 52.890 31.040 53.290 32.140 ;
        RECT 54.890 31.040 55.290 32.140 ;
        RECT 56.890 31.040 57.290 32.140 ;
        RECT 58.890 31.040 59.290 32.140 ;
        RECT 60.890 31.040 61.290 32.140 ;
        RECT 62.890 31.040 63.290 32.140 ;
        RECT 64.890 31.040 65.290 32.140 ;
        RECT 66.890 31.040 67.290 32.140 ;
        RECT 68.890 31.040 69.290 32.140 ;
        RECT 70.890 31.040 71.290 32.140 ;
        RECT 72.890 31.040 73.290 32.140 ;
        RECT 6.890 29.190 7.290 30.290 ;
        RECT 8.890 29.190 9.290 30.290 ;
        RECT 10.890 29.190 11.290 30.290 ;
        RECT 12.890 29.190 13.290 30.290 ;
        RECT 14.890 29.190 15.290 30.290 ;
        RECT 16.890 29.190 17.290 30.290 ;
        RECT 18.890 29.190 19.290 30.290 ;
        RECT 20.890 29.190 21.290 30.290 ;
        RECT 22.890 29.190 23.290 30.290 ;
        RECT 24.890 29.190 25.290 30.290 ;
        RECT 26.890 29.190 27.290 30.290 ;
        RECT 28.890 29.190 29.290 30.290 ;
        RECT 30.890 29.190 31.290 30.290 ;
        RECT 32.890 29.190 33.290 30.290 ;
        RECT 34.890 29.190 35.290 30.290 ;
        RECT 36.890 29.190 37.290 30.290 ;
        RECT 38.890 29.190 39.290 30.290 ;
        RECT 40.890 29.190 41.290 30.290 ;
        RECT 42.890 29.190 43.290 30.290 ;
        RECT 44.890 29.190 45.290 30.290 ;
        RECT 46.890 29.190 47.290 30.290 ;
        RECT 48.890 29.190 49.290 30.290 ;
        RECT 50.890 29.190 51.290 30.290 ;
        RECT 52.890 29.190 53.290 30.290 ;
        RECT 54.890 29.190 55.290 30.290 ;
        RECT 56.890 29.190 57.290 30.290 ;
        RECT 58.890 29.190 59.290 30.290 ;
        RECT 60.890 29.190 61.290 30.290 ;
        RECT 62.890 29.190 63.290 30.290 ;
        RECT 64.890 29.190 65.290 30.290 ;
        RECT 66.890 29.190 67.290 30.290 ;
        RECT 68.890 29.190 69.290 30.290 ;
        RECT 70.890 29.190 71.290 30.290 ;
        RECT 72.890 29.190 73.290 30.290 ;
        RECT 6.890 27.340 7.290 28.440 ;
        RECT 8.890 27.340 9.290 28.440 ;
        RECT 10.890 27.340 11.290 28.440 ;
        RECT 12.890 27.340 13.290 28.440 ;
        RECT 14.890 27.340 15.290 28.440 ;
        RECT 16.890 27.340 17.290 28.440 ;
        RECT 18.890 27.340 19.290 28.440 ;
        RECT 20.890 27.340 21.290 28.440 ;
        RECT 22.890 27.340 23.290 28.440 ;
        RECT 24.890 27.340 25.290 28.440 ;
        RECT 26.890 27.340 27.290 28.440 ;
        RECT 28.890 27.340 29.290 28.440 ;
        RECT 30.890 27.340 31.290 28.440 ;
        RECT 32.890 27.340 33.290 28.440 ;
        RECT 34.890 27.340 35.290 28.440 ;
        RECT 36.890 27.340 37.290 28.440 ;
        RECT 38.890 27.340 39.290 28.440 ;
        RECT 40.890 27.340 41.290 28.440 ;
        RECT 42.890 27.340 43.290 28.440 ;
        RECT 44.890 27.340 45.290 28.440 ;
        RECT 46.890 27.340 47.290 28.440 ;
        RECT 48.890 27.340 49.290 28.440 ;
        RECT 50.890 27.340 51.290 28.440 ;
        RECT 52.890 27.340 53.290 28.440 ;
        RECT 54.890 27.340 55.290 28.440 ;
        RECT 56.890 27.340 57.290 28.440 ;
        RECT 58.890 27.340 59.290 28.440 ;
        RECT 60.890 27.340 61.290 28.440 ;
        RECT 62.890 27.340 63.290 28.440 ;
        RECT 64.890 27.340 65.290 28.440 ;
        RECT 66.890 27.340 67.290 28.440 ;
        RECT 68.890 27.340 69.290 28.440 ;
        RECT 70.890 27.340 71.290 28.440 ;
        RECT 72.890 27.340 73.290 28.440 ;
        RECT 6.890 25.490 7.290 26.590 ;
        RECT 8.890 25.490 9.290 26.590 ;
        RECT 10.890 25.490 11.290 26.590 ;
        RECT 12.890 25.490 13.290 26.590 ;
        RECT 14.890 25.490 15.290 26.590 ;
        RECT 16.890 25.490 17.290 26.590 ;
        RECT 18.890 25.490 19.290 26.590 ;
        RECT 20.890 25.490 21.290 26.590 ;
        RECT 22.890 25.490 23.290 26.590 ;
        RECT 24.890 25.490 25.290 26.590 ;
        RECT 26.890 25.490 27.290 26.590 ;
        RECT 28.890 25.490 29.290 26.590 ;
        RECT 30.890 25.490 31.290 26.590 ;
        RECT 32.890 25.490 33.290 26.590 ;
        RECT 34.890 25.490 35.290 26.590 ;
        RECT 36.890 25.490 37.290 26.590 ;
        RECT 38.890 25.490 39.290 26.590 ;
        RECT 40.890 25.490 41.290 26.590 ;
        RECT 42.890 25.490 43.290 26.590 ;
        RECT 44.890 25.490 45.290 26.590 ;
        RECT 46.890 25.490 47.290 26.590 ;
        RECT 48.890 25.490 49.290 26.590 ;
        RECT 50.890 25.490 51.290 26.590 ;
        RECT 52.890 25.490 53.290 26.590 ;
        RECT 54.890 25.490 55.290 26.590 ;
        RECT 56.890 25.490 57.290 26.590 ;
        RECT 58.890 25.490 59.290 26.590 ;
        RECT 60.890 25.490 61.290 26.590 ;
        RECT 62.890 25.490 63.290 26.590 ;
        RECT 64.890 25.490 65.290 26.590 ;
        RECT 66.890 25.490 67.290 26.590 ;
        RECT 68.890 25.490 69.290 26.590 ;
        RECT 70.890 25.490 71.290 26.590 ;
        RECT 72.890 25.490 73.290 26.590 ;
        RECT 75.040 26.240 75.240 132.340 ;
        RECT 75.440 131.890 75.740 132.290 ;
        RECT 85.375 131.890 85.675 132.290 ;
        RECT 75.490 37.340 75.690 131.890 ;
        RECT 75.890 131.440 76.190 131.840 ;
        RECT 84.925 131.440 85.225 131.840 ;
        RECT 75.940 46.590 76.140 131.440 ;
        RECT 76.340 130.990 76.640 131.390 ;
        RECT 84.475 130.990 84.775 131.390 ;
        RECT 76.390 52.140 76.590 130.990 ;
        RECT 76.790 130.540 77.090 130.940 ;
        RECT 84.025 130.540 84.325 130.940 ;
        RECT 76.840 55.840 77.040 130.540 ;
        RECT 77.240 130.090 77.540 130.490 ;
        RECT 83.575 130.090 83.875 130.490 ;
        RECT 77.290 57.690 77.490 130.090 ;
        RECT 77.690 129.640 77.990 130.040 ;
        RECT 83.125 129.640 83.425 130.040 ;
        RECT 77.740 61.390 77.940 129.640 ;
        RECT 79.940 129.190 80.240 129.590 ;
        RECT 80.875 129.190 81.175 129.590 ;
        RECT 78.140 128.740 78.440 129.140 ;
        RECT 78.190 63.240 78.390 128.740 ;
        RECT 79.490 128.290 79.790 128.690 ;
        RECT 79.040 127.840 79.340 128.240 ;
        RECT 78.590 127.390 78.890 127.790 ;
        RECT 78.640 65.090 78.840 127.390 ;
        RECT 79.090 66.940 79.290 127.840 ;
        RECT 79.540 68.790 79.740 128.290 ;
        RECT 79.990 70.640 80.190 129.190 ;
        RECT 80.925 70.640 81.125 129.190 ;
        RECT 82.675 128.740 82.975 129.140 ;
        RECT 81.325 128.290 81.625 128.690 ;
        RECT 79.940 70.240 80.240 70.640 ;
        RECT 80.875 70.240 81.175 70.640 ;
        RECT 81.375 68.790 81.575 128.290 ;
        RECT 81.775 127.840 82.075 128.240 ;
        RECT 79.490 68.390 79.790 68.790 ;
        RECT 81.325 68.390 81.625 68.790 ;
        RECT 81.825 66.940 82.025 127.840 ;
        RECT 82.225 127.390 82.525 127.790 ;
        RECT 79.040 66.540 79.340 66.940 ;
        RECT 81.775 66.540 82.075 66.940 ;
        RECT 82.275 65.090 82.475 127.390 ;
        RECT 78.590 64.690 78.890 65.090 ;
        RECT 82.225 64.690 82.525 65.090 ;
        RECT 82.725 63.240 82.925 128.740 ;
        RECT 78.140 62.840 78.440 63.240 ;
        RECT 82.675 62.840 82.975 63.240 ;
        RECT 83.175 61.390 83.375 129.640 ;
        RECT 77.690 60.990 77.990 61.390 ;
        RECT 83.125 60.990 83.425 61.390 ;
        RECT 83.625 57.690 83.825 130.090 ;
        RECT 77.240 57.290 77.540 57.690 ;
        RECT 83.575 57.290 83.875 57.690 ;
        RECT 84.075 55.840 84.275 130.540 ;
        RECT 76.790 55.440 77.090 55.840 ;
        RECT 84.025 55.440 84.325 55.840 ;
        RECT 84.525 52.140 84.725 130.990 ;
        RECT 76.340 51.740 76.640 52.140 ;
        RECT 84.475 51.740 84.775 52.140 ;
        RECT 84.975 46.590 85.175 131.440 ;
        RECT 75.890 46.190 76.190 46.590 ;
        RECT 84.925 46.190 85.225 46.590 ;
        RECT 85.425 37.340 85.625 131.890 ;
        RECT 75.440 36.940 75.740 37.340 ;
        RECT 85.375 36.940 85.675 37.340 ;
        RECT 85.875 26.240 86.075 132.340 ;
        RECT 86.375 127.790 86.575 141.015 ;
        RECT 88.225 139.565 88.375 141.215 ;
        RECT 86.725 139.015 87.025 139.415 ;
        RECT 88.125 139.165 88.425 139.565 ;
        RECT 92.725 139.215 92.925 143.290 ;
        RECT 86.775 128.690 86.975 139.015 ;
        RECT 88.225 137.415 88.375 139.165 ;
        RECT 92.675 138.815 92.975 139.215 ;
        RECT 93.125 138.015 93.325 145.090 ;
        RECT 93.475 143.740 93.775 144.140 ;
        RECT 93.525 138.815 93.725 143.740 ;
        RECT 93.475 138.415 93.775 138.815 ;
        RECT 93.075 137.615 93.375 138.015 ;
        RECT 93.925 137.615 94.125 145.540 ;
        RECT 94.275 144.190 94.575 144.590 ;
        RECT 94.325 138.415 94.525 144.190 ;
        RECT 94.275 138.015 94.575 138.415 ;
        RECT 87.125 136.765 87.425 137.165 ;
        RECT 88.125 137.015 88.425 137.415 ;
        RECT 93.875 137.215 94.175 137.615 ;
        RECT 94.725 137.215 94.925 145.990 ;
        RECT 95.075 144.640 95.375 145.040 ;
        RECT 87.175 129.590 87.375 136.765 ;
        RECT 87.575 135.615 87.875 135.715 ;
        RECT 88.225 135.615 88.375 137.015 ;
        RECT 94.675 136.815 94.975 137.215 ;
        RECT 95.125 136.265 95.325 144.640 ;
        RECT 95.525 136.815 95.725 146.440 ;
        RECT 101.875 145.990 102.175 146.390 ;
        RECT 100.925 145.540 101.225 145.940 ;
        RECT 100.325 145.090 100.625 145.490 ;
        RECT 99.275 144.640 99.575 145.040 ;
        RECT 98.225 144.190 98.525 144.590 ;
        RECT 97.175 143.740 97.475 144.140 ;
        RECT 96.125 143.290 96.425 143.690 ;
        RECT 96.175 142.265 96.375 143.290 ;
        RECT 97.225 142.265 97.425 143.740 ;
        RECT 98.275 142.265 98.475 144.190 ;
        RECT 99.325 142.265 99.525 144.640 ;
        RECT 100.375 142.265 100.575 145.090 ;
        RECT 100.975 142.265 101.175 145.540 ;
        RECT 101.925 142.265 102.125 145.990 ;
        RECT 102.975 142.265 103.175 146.890 ;
        RECT 103.925 142.265 104.125 147.340 ;
        RECT 105.825 142.265 106.025 147.790 ;
        RECT 109.675 142.265 109.875 148.240 ;
        RECT 113.525 142.265 113.725 148.690 ;
        RECT 123.325 148.240 123.625 148.640 ;
        RECT 119.475 147.790 119.775 148.190 ;
        RECT 117.525 147.340 117.825 147.740 ;
        RECT 116.675 146.890 116.975 147.290 ;
        RECT 115.575 146.440 115.875 146.840 ;
        RECT 115.625 142.265 115.825 146.440 ;
        RECT 116.725 142.265 116.925 146.890 ;
        RECT 117.575 142.265 117.775 147.340 ;
        RECT 119.525 142.265 119.725 147.790 ;
        RECT 123.375 142.265 123.575 148.240 ;
        RECT 124.275 146.840 124.475 152.890 ;
        RECT 127.540 152.590 129.390 153.690 ;
        RECT 150.850 153.490 151.250 153.540 ;
        RECT 155.525 153.490 155.875 153.690 ;
        RECT 150.850 153.290 152.775 153.490 ;
        RECT 150.850 153.240 151.250 153.290 ;
        RECT 142.250 152.740 142.550 153.140 ;
        RECT 137.175 152.290 137.475 152.690 ;
        RECT 134.575 151.840 134.875 152.240 ;
        RECT 133.325 151.390 133.625 151.790 ;
        RECT 132.125 150.940 132.425 151.340 ;
        RECT 130.875 150.490 131.175 150.890 ;
        RECT 129.675 150.040 129.975 150.440 ;
        RECT 128.475 149.590 128.775 149.990 ;
        RECT 127.225 149.140 127.525 149.540 ;
        RECT 126.075 148.690 126.375 149.090 ;
        RECT 124.225 146.440 124.525 146.840 ;
        RECT 126.125 142.365 126.325 148.690 ;
        RECT 127.275 142.365 127.475 149.140 ;
        RECT 128.525 142.365 128.725 149.590 ;
        RECT 129.725 142.365 129.925 150.040 ;
        RECT 130.925 142.365 131.125 150.490 ;
        RECT 132.175 142.365 132.375 150.940 ;
        RECT 133.375 142.365 133.575 151.390 ;
        RECT 134.625 142.365 134.825 151.840 ;
        RECT 137.225 142.365 137.425 152.290 ;
        RECT 142.350 143.565 142.550 152.740 ;
        RECT 142.300 143.140 142.550 143.565 ;
        RECT 142.300 142.365 142.500 143.140 ;
        RECT 152.575 142.365 152.775 153.290 ;
        RECT 96.125 141.865 96.425 142.265 ;
        RECT 97.175 141.865 97.475 142.265 ;
        RECT 98.225 141.865 98.525 142.265 ;
        RECT 99.275 141.865 99.575 142.265 ;
        RECT 100.325 141.865 100.625 142.265 ;
        RECT 100.925 141.865 101.225 142.265 ;
        RECT 101.875 141.865 102.175 142.265 ;
        RECT 102.925 141.865 103.225 142.265 ;
        RECT 103.875 141.865 104.175 142.265 ;
        RECT 105.775 141.865 106.075 142.265 ;
        RECT 109.625 141.865 109.925 142.265 ;
        RECT 113.475 141.865 113.775 142.265 ;
        RECT 115.575 141.865 115.875 142.265 ;
        RECT 116.675 141.865 116.975 142.265 ;
        RECT 117.525 141.865 117.825 142.265 ;
        RECT 119.475 141.865 119.775 142.265 ;
        RECT 123.325 141.865 123.625 142.265 ;
        RECT 126.075 141.965 126.375 142.365 ;
        RECT 127.225 141.965 127.525 142.365 ;
        RECT 128.475 141.965 128.775 142.365 ;
        RECT 129.675 141.965 129.975 142.365 ;
        RECT 130.875 141.965 131.175 142.365 ;
        RECT 132.125 141.965 132.425 142.365 ;
        RECT 133.325 141.965 133.625 142.365 ;
        RECT 134.575 141.965 134.875 142.365 ;
        RECT 137.175 141.965 137.475 142.365 ;
        RECT 142.275 141.965 142.575 142.365 ;
        RECT 152.475 141.965 152.875 142.365 ;
        RECT 103.625 141.565 103.925 141.665 ;
        RECT 104.575 141.565 104.875 141.665 ;
        RECT 105.525 141.565 105.825 141.665 ;
        RECT 106.475 141.565 106.775 141.665 ;
        RECT 107.475 141.565 107.775 141.665 ;
        RECT 108.425 141.565 108.725 141.665 ;
        RECT 109.375 141.565 109.675 141.665 ;
        RECT 110.325 141.565 110.625 141.665 ;
        RECT 111.325 141.565 111.625 141.665 ;
        RECT 112.275 141.565 112.575 141.665 ;
        RECT 113.225 141.565 113.525 141.665 ;
        RECT 114.175 141.565 114.475 141.665 ;
        RECT 154.925 141.565 155.225 141.640 ;
        RECT 103.625 141.365 155.225 141.565 ;
        RECT 103.625 141.265 103.925 141.365 ;
        RECT 104.575 141.215 104.875 141.365 ;
        RECT 105.525 141.265 105.825 141.365 ;
        RECT 106.475 141.265 106.775 141.365 ;
        RECT 107.475 141.265 107.775 141.365 ;
        RECT 108.425 141.265 108.725 141.365 ;
        RECT 109.375 141.265 109.675 141.365 ;
        RECT 110.325 141.265 110.625 141.365 ;
        RECT 111.325 141.265 111.625 141.365 ;
        RECT 112.275 141.265 112.575 141.365 ;
        RECT 113.225 141.265 113.525 141.365 ;
        RECT 114.175 141.265 114.475 141.365 ;
        RECT 154.925 141.240 155.225 141.365 ;
        RECT 96.375 141.065 96.675 141.165 ;
        RECT 97.425 141.065 97.725 141.165 ;
        RECT 98.475 141.065 98.775 141.165 ;
        RECT 99.525 141.065 99.825 141.165 ;
        RECT 100.575 141.065 100.875 141.165 ;
        RECT 101.625 141.065 101.925 141.165 ;
        RECT 102.575 141.065 102.875 141.165 ;
        RECT 96.375 140.865 103.925 141.065 ;
        RECT 96.375 140.765 96.675 140.865 ;
        RECT 97.425 140.765 97.725 140.865 ;
        RECT 98.475 140.765 98.775 140.865 ;
        RECT 99.525 140.765 99.825 140.865 ;
        RECT 100.575 140.765 100.875 140.865 ;
        RECT 101.625 140.765 101.925 140.865 ;
        RECT 102.575 140.815 103.925 140.865 ;
        RECT 102.575 140.765 102.825 140.815 ;
        RECT 103.625 140.665 103.925 140.815 ;
        RECT 110.825 140.565 111.125 140.665 ;
        RECT 111.775 140.565 112.075 140.665 ;
        RECT 112.225 140.565 112.525 140.665 ;
        RECT 112.725 140.565 113.025 140.665 ;
        RECT 113.675 140.565 113.975 140.665 ;
        RECT 110.825 140.365 113.975 140.565 ;
        RECT 95.875 139.965 96.175 140.365 ;
        RECT 96.925 139.965 97.225 140.365 ;
        RECT 97.975 139.915 98.275 140.315 ;
        RECT 99.025 139.915 99.325 140.315 ;
        RECT 100.075 139.915 100.375 140.315 ;
        RECT 101.125 139.915 101.425 140.315 ;
        RECT 102.075 139.915 102.375 140.315 ;
        RECT 110.825 140.265 111.125 140.365 ;
        RECT 111.775 140.265 112.075 140.365 ;
        RECT 112.225 140.265 112.525 140.365 ;
        RECT 112.725 140.265 113.025 140.365 ;
        RECT 113.675 140.265 113.975 140.365 ;
        RECT 96.625 139.515 96.925 139.615 ;
        RECT 115.575 139.515 115.875 139.615 ;
        RECT 96.625 139.315 115.875 139.515 ;
        RECT 96.625 139.215 96.925 139.315 ;
        RECT 115.575 139.215 115.875 139.315 ;
        RECT 100.875 138.415 101.175 138.815 ;
        RECT 101.825 138.765 102.125 139.165 ;
        RECT 100.325 138.015 100.625 138.415 ;
        RECT 99.275 137.615 99.575 138.015 ;
        RECT 98.225 137.215 98.525 137.615 ;
        RECT 97.175 136.815 97.475 137.215 ;
        RECT 95.475 136.415 95.775 136.815 ;
        RECT 96.125 136.415 96.425 136.815 ;
        RECT 96.175 136.265 96.375 136.415 ;
        RECT 97.225 136.265 97.425 136.815 ;
        RECT 98.275 136.265 98.475 137.215 ;
        RECT 99.325 136.265 99.525 137.615 ;
        RECT 100.375 136.265 100.575 138.015 ;
        RECT 100.925 136.265 101.125 138.415 ;
        RECT 101.875 136.265 102.075 138.765 ;
        RECT 103.625 138.365 103.925 138.465 ;
        RECT 117.325 138.365 117.625 138.465 ;
        RECT 103.625 138.165 117.625 138.365 ;
        RECT 124.040 138.240 125.840 140.140 ;
        RECT 153.475 140.065 153.775 140.915 ;
        RECT 155.575 140.065 155.875 140.140 ;
        RECT 153.475 139.865 155.875 140.065 ;
        RECT 153.475 139.015 153.775 139.865 ;
        RECT 155.575 139.740 155.875 139.865 ;
        RECT 126.375 138.515 126.675 138.615 ;
        RECT 127.575 138.515 127.875 138.615 ;
        RECT 128.775 138.515 129.075 138.615 ;
        RECT 130.025 138.515 130.325 138.615 ;
        RECT 131.225 138.515 131.525 138.615 ;
        RECT 132.425 138.515 132.725 138.615 ;
        RECT 133.625 138.515 133.925 138.615 ;
        RECT 134.925 138.515 135.225 138.615 ;
        RECT 136.225 138.515 136.525 138.615 ;
        RECT 137.475 138.515 137.775 138.615 ;
        RECT 138.775 138.515 139.075 138.615 ;
        RECT 140.075 138.515 140.375 138.615 ;
        RECT 141.325 138.515 141.625 138.615 ;
        RECT 142.625 138.515 142.925 138.615 ;
        RECT 143.875 138.515 144.175 138.615 ;
        RECT 145.175 138.515 145.475 138.615 ;
        RECT 146.475 138.515 146.775 138.615 ;
        RECT 147.725 138.515 148.025 138.615 ;
        RECT 149.025 138.515 149.325 138.615 ;
        RECT 150.275 138.515 150.575 138.615 ;
        RECT 151.575 138.515 151.875 138.615 ;
        RECT 152.875 138.515 153.175 138.615 ;
        RECT 156.225 138.515 156.525 138.590 ;
        RECT 126.375 138.315 156.525 138.515 ;
        RECT 126.375 138.215 126.675 138.315 ;
        RECT 127.575 138.215 127.875 138.315 ;
        RECT 128.775 138.215 129.075 138.315 ;
        RECT 130.025 138.215 130.325 138.315 ;
        RECT 131.225 138.215 131.525 138.315 ;
        RECT 132.425 138.215 132.725 138.315 ;
        RECT 133.625 138.215 133.925 138.315 ;
        RECT 134.925 138.215 135.225 138.315 ;
        RECT 136.225 138.215 136.525 138.315 ;
        RECT 137.475 138.215 137.775 138.315 ;
        RECT 138.775 138.215 139.075 138.315 ;
        RECT 140.075 138.215 140.375 138.315 ;
        RECT 141.325 138.215 141.625 138.315 ;
        RECT 142.625 138.215 142.925 138.315 ;
        RECT 143.875 138.215 144.175 138.315 ;
        RECT 145.175 138.215 145.475 138.315 ;
        RECT 146.475 138.215 146.775 138.315 ;
        RECT 147.725 138.215 148.025 138.315 ;
        RECT 149.025 138.215 149.325 138.315 ;
        RECT 150.275 138.215 150.575 138.315 ;
        RECT 151.575 138.215 151.875 138.315 ;
        RECT 152.875 138.215 153.175 138.315 ;
        RECT 156.225 138.190 156.525 138.315 ;
        RECT 103.625 138.065 103.925 138.165 ;
        RECT 117.325 138.065 117.625 138.165 ;
        RECT 117.325 136.465 117.625 136.565 ;
        RECT 118.275 136.465 118.575 136.565 ;
        RECT 119.225 136.465 119.525 136.565 ;
        RECT 120.175 136.465 120.475 136.565 ;
        RECT 121.125 136.465 121.425 136.565 ;
        RECT 122.125 136.465 122.425 136.565 ;
        RECT 123.075 136.465 123.375 136.565 ;
        RECT 124.025 136.465 124.325 136.565 ;
        RECT 156.875 136.465 157.175 136.540 ;
        RECT 117.325 136.265 157.175 136.465 ;
        RECT 95.075 135.865 95.375 136.265 ;
        RECT 96.125 135.865 96.425 136.265 ;
        RECT 97.175 135.865 97.475 136.265 ;
        RECT 98.225 135.865 98.525 136.265 ;
        RECT 99.275 135.865 99.575 136.265 ;
        RECT 100.325 135.865 100.625 136.265 ;
        RECT 100.875 135.865 101.175 136.265 ;
        RECT 101.825 135.865 102.125 136.265 ;
        RECT 117.325 136.165 117.625 136.265 ;
        RECT 118.275 136.165 118.575 136.265 ;
        RECT 119.225 136.165 119.525 136.265 ;
        RECT 120.175 136.165 120.475 136.265 ;
        RECT 121.125 136.165 121.425 136.265 ;
        RECT 122.125 136.165 122.425 136.265 ;
        RECT 123.075 136.165 123.375 136.265 ;
        RECT 124.025 136.165 124.325 136.265 ;
        RECT 156.875 136.140 157.175 136.265 ;
        RECT 115.325 135.815 115.625 135.915 ;
        RECT 116.275 135.815 116.575 135.915 ;
        RECT 157.525 135.815 157.825 135.890 ;
        RECT 88.625 135.615 88.925 135.715 ;
        RECT 89.675 135.615 89.975 135.715 ;
        RECT 90.725 135.615 91.025 135.715 ;
        RECT 91.775 135.615 92.075 135.715 ;
        RECT 93.325 135.615 93.625 135.715 ;
        RECT 94.275 135.615 94.575 135.715 ;
        RECT 87.575 135.415 94.575 135.615 ;
        RECT 87.575 135.315 87.875 135.415 ;
        RECT 88.625 135.315 88.925 135.415 ;
        RECT 89.675 135.315 89.975 135.415 ;
        RECT 90.725 135.315 91.025 135.415 ;
        RECT 91.775 135.315 92.075 135.415 ;
        RECT 93.325 135.315 93.625 135.415 ;
        RECT 94.275 135.315 94.575 135.415 ;
        RECT 95.325 135.665 95.625 135.715 ;
        RECT 96.375 135.665 96.675 135.715 ;
        RECT 97.425 135.665 97.725 135.715 ;
        RECT 98.475 135.665 98.775 135.715 ;
        RECT 99.525 135.665 99.825 135.715 ;
        RECT 100.575 135.665 100.875 135.715 ;
        RECT 101.625 135.665 101.925 135.715 ;
        RECT 102.575 135.665 102.875 135.715 ;
        RECT 104.575 135.665 104.875 135.715 ;
        RECT 95.325 135.365 104.875 135.665 ;
        RECT 115.325 135.615 157.825 135.815 ;
        RECT 115.325 135.515 115.650 135.615 ;
        RECT 116.275 135.515 116.575 135.615 ;
        RECT 95.325 135.315 95.625 135.365 ;
        RECT 96.375 135.315 96.675 135.365 ;
        RECT 97.425 135.315 97.725 135.365 ;
        RECT 98.475 135.315 98.775 135.365 ;
        RECT 99.525 135.315 99.825 135.365 ;
        RECT 100.575 135.315 100.875 135.365 ;
        RECT 101.625 135.315 101.925 135.365 ;
        RECT 102.575 135.315 102.875 135.365 ;
        RECT 104.575 135.315 104.875 135.365 ;
        RECT 88.075 134.765 88.375 135.165 ;
        RECT 89.125 134.765 89.425 135.165 ;
        RECT 90.175 134.765 90.475 135.165 ;
        RECT 91.225 134.765 91.525 135.165 ;
        RECT 92.275 134.765 92.575 135.165 ;
        RECT 94.325 134.965 94.475 135.315 ;
        RECT 115.400 134.965 115.650 135.515 ;
        RECT 157.525 135.490 157.825 135.615 ;
        RECT 87.125 129.190 87.425 129.590 ;
        RECT 86.725 128.290 87.025 128.690 ;
        RECT 88.125 128.240 88.325 134.765 ;
        RECT 89.175 129.140 89.375 134.765 ;
        RECT 90.225 130.040 90.425 134.765 ;
        RECT 91.275 130.490 91.475 134.765 ;
        RECT 92.325 130.940 92.525 134.765 ;
        RECT 94.325 134.715 115.650 134.965 ;
        RECT 92.825 133.865 93.125 134.265 ;
        RECT 93.775 133.865 94.075 134.265 ;
        RECT 94.825 134.015 95.125 134.415 ;
        RECT 95.875 134.015 96.175 134.415 ;
        RECT 96.925 134.015 97.225 134.415 ;
        RECT 97.975 134.015 98.275 134.415 ;
        RECT 99.025 134.015 99.325 134.415 ;
        RECT 100.075 134.015 100.375 134.415 ;
        RECT 101.125 134.015 101.425 134.415 ;
        RECT 102.075 134.015 102.375 134.415 ;
        RECT 92.875 131.390 93.075 133.865 ;
        RECT 93.825 131.840 94.025 133.865 ;
        RECT 93.775 131.440 94.075 131.840 ;
        RECT 92.825 130.990 93.125 131.390 ;
        RECT 92.275 130.540 92.575 130.940 ;
        RECT 91.225 130.090 91.525 130.490 ;
        RECT 90.175 129.640 90.475 130.040 ;
        RECT 89.125 128.740 89.425 129.140 ;
        RECT 88.075 127.840 88.375 128.240 ;
        RECT 94.875 127.790 95.075 134.015 ;
        RECT 95.925 128.240 96.125 134.015 ;
        RECT 96.975 128.690 97.175 134.015 ;
        RECT 98.025 129.140 98.225 134.015 ;
        RECT 99.075 129.590 99.275 134.015 ;
        RECT 100.125 130.040 100.325 134.015 ;
        RECT 101.175 130.490 101.375 134.015 ;
        RECT 102.125 130.940 102.325 134.015 ;
        RECT 103.125 133.815 103.425 134.215 ;
        RECT 104.075 133.815 104.375 134.215 ;
        RECT 105.075 134.115 105.375 134.215 ;
        RECT 106.025 134.115 106.325 134.215 ;
        RECT 105.075 133.915 106.325 134.115 ;
        RECT 105.075 133.815 105.375 133.915 ;
        RECT 106.025 133.815 106.325 133.915 ;
        RECT 106.975 134.115 107.275 134.215 ;
        RECT 107.925 134.115 108.225 134.215 ;
        RECT 108.875 134.115 109.175 134.215 ;
        RECT 109.875 134.115 110.175 134.215 ;
        RECT 106.975 133.915 110.175 134.115 ;
        RECT 114.825 133.965 115.125 134.365 ;
        RECT 115.775 133.965 116.075 134.365 ;
        RECT 116.825 133.965 117.125 134.365 ;
        RECT 117.775 133.965 118.075 134.365 ;
        RECT 118.725 134.265 119.025 134.365 ;
        RECT 119.725 134.265 120.025 134.365 ;
        RECT 118.725 134.065 120.025 134.265 ;
        RECT 118.725 133.965 119.025 134.065 ;
        RECT 119.725 133.965 120.025 134.065 ;
        RECT 120.675 134.265 120.975 134.365 ;
        RECT 121.625 134.265 121.925 134.365 ;
        RECT 122.575 134.265 122.875 134.365 ;
        RECT 123.525 134.265 123.825 134.365 ;
        RECT 120.675 134.065 123.825 134.265 ;
        RECT 120.675 133.965 120.975 134.065 ;
        RECT 121.625 133.965 121.925 134.065 ;
        RECT 122.575 133.965 122.875 134.065 ;
        RECT 123.525 133.965 123.825 134.065 ;
        RECT 106.975 133.815 107.275 133.915 ;
        RECT 107.925 133.815 108.225 133.915 ;
        RECT 108.875 133.815 109.175 133.915 ;
        RECT 109.875 133.815 110.175 133.915 ;
        RECT 103.175 131.390 103.375 133.815 ;
        RECT 104.175 131.840 104.375 133.815 ;
        RECT 106.075 132.290 106.275 133.815 ;
        RECT 106.675 133.040 109.525 133.440 ;
        RECT 109.925 132.740 110.125 133.815 ;
        RECT 109.875 132.340 110.175 132.740 ;
        RECT 114.875 132.290 115.075 133.965 ;
        RECT 115.825 132.740 116.025 133.965 ;
        RECT 115.775 132.340 116.075 132.740 ;
        RECT 106.025 131.890 106.325 132.290 ;
        RECT 114.825 131.890 115.125 132.290 ;
        RECT 104.125 131.440 104.425 131.840 ;
        RECT 116.875 131.390 117.075 133.965 ;
        RECT 117.825 131.840 118.025 133.965 ;
        RECT 119.775 132.290 119.975 133.965 ;
        RECT 120.325 133.040 123.175 133.440 ;
        RECT 123.575 132.740 123.775 133.965 ;
        RECT 125.725 133.715 126.025 134.115 ;
        RECT 126.925 133.715 127.225 134.115 ;
        RECT 128.125 133.715 128.425 134.115 ;
        RECT 129.375 133.715 129.675 134.115 ;
        RECT 130.575 133.715 130.875 134.115 ;
        RECT 131.775 133.715 132.075 134.115 ;
        RECT 133.025 133.865 133.325 134.265 ;
        RECT 134.275 133.865 134.575 134.265 ;
        RECT 135.575 134.165 135.875 134.265 ;
        RECT 136.875 134.165 137.175 134.265 ;
        RECT 135.575 133.965 137.175 134.165 ;
        RECT 135.575 133.865 135.875 133.965 ;
        RECT 136.875 133.865 137.175 133.965 ;
        RECT 138.125 134.165 138.425 134.265 ;
        RECT 139.425 134.165 139.725 134.265 ;
        RECT 140.675 134.165 140.975 134.265 ;
        RECT 141.975 134.165 142.275 134.265 ;
        RECT 138.125 133.965 142.275 134.165 ;
        RECT 138.125 133.865 138.425 133.965 ;
        RECT 139.425 133.865 139.725 133.965 ;
        RECT 140.675 133.865 140.975 133.965 ;
        RECT 141.975 133.865 142.275 133.965 ;
        RECT 143.225 134.165 143.525 134.265 ;
        RECT 144.525 134.165 144.825 134.265 ;
        RECT 145.825 134.165 146.125 134.265 ;
        RECT 147.075 134.165 147.375 134.265 ;
        RECT 148.375 134.165 148.675 134.265 ;
        RECT 149.625 134.165 149.925 134.265 ;
        RECT 150.925 134.165 151.225 134.265 ;
        RECT 152.225 134.165 152.525 134.265 ;
        RECT 143.225 133.965 152.525 134.165 ;
        RECT 143.225 133.865 143.525 133.965 ;
        RECT 144.525 133.865 144.825 133.965 ;
        RECT 145.825 133.865 146.125 133.965 ;
        RECT 147.075 133.865 147.375 133.965 ;
        RECT 148.375 133.865 148.675 133.965 ;
        RECT 149.625 133.865 149.925 133.965 ;
        RECT 150.925 133.865 151.225 133.965 ;
        RECT 152.225 133.865 152.525 133.965 ;
        RECT 123.525 132.340 123.825 132.740 ;
        RECT 119.725 131.890 120.025 132.290 ;
        RECT 117.775 131.440 118.075 131.840 ;
        RECT 103.125 130.990 103.425 131.390 ;
        RECT 116.825 130.990 117.125 131.390 ;
        RECT 102.075 130.540 102.375 130.940 ;
        RECT 101.125 130.090 101.425 130.490 ;
        RECT 100.075 129.640 100.375 130.040 ;
        RECT 99.025 129.190 99.325 129.590 ;
        RECT 97.975 128.740 98.275 129.140 ;
        RECT 96.925 128.290 97.225 128.690 ;
        RECT 125.775 128.240 125.975 133.715 ;
        RECT 126.975 128.690 127.175 133.715 ;
        RECT 128.175 129.140 128.375 133.715 ;
        RECT 129.425 129.590 129.625 133.715 ;
        RECT 130.625 130.040 130.825 133.715 ;
        RECT 131.825 130.490 132.025 133.715 ;
        RECT 133.075 130.940 133.275 133.865 ;
        RECT 134.325 131.390 134.525 133.865 ;
        RECT 136.925 131.840 137.125 133.865 ;
        RECT 142.025 132.290 142.225 133.865 ;
        RECT 152.275 132.740 152.475 133.865 ;
        RECT 152.225 132.340 152.525 132.740 ;
        RECT 141.975 131.890 142.275 132.290 ;
        RECT 136.875 131.440 137.175 131.840 ;
        RECT 134.275 130.990 134.575 131.390 ;
        RECT 133.025 130.540 133.325 130.940 ;
        RECT 131.775 130.090 132.075 130.490 ;
        RECT 130.575 129.640 130.875 130.040 ;
        RECT 129.375 129.190 129.675 129.590 ;
        RECT 128.125 128.740 128.425 129.140 ;
        RECT 126.925 128.290 127.225 128.690 ;
        RECT 95.875 127.840 96.175 128.240 ;
        RECT 125.725 127.840 126.025 128.240 ;
        RECT 86.325 127.390 86.625 127.790 ;
        RECT 94.825 127.390 95.125 127.790 ;
        RECT 86.825 126.940 87.725 127.340 ;
        RECT 152.825 127.190 153.725 127.590 ;
        RECT 87.825 125.390 88.225 126.490 ;
        RECT 89.825 125.390 90.225 126.490 ;
        RECT 91.825 125.390 92.225 126.490 ;
        RECT 93.825 125.390 94.225 126.490 ;
        RECT 95.825 125.390 96.225 126.490 ;
        RECT 97.825 125.390 98.225 126.490 ;
        RECT 99.825 125.390 100.225 126.490 ;
        RECT 101.825 125.390 102.225 126.490 ;
        RECT 103.825 125.390 104.225 126.490 ;
        RECT 105.825 125.390 106.225 126.490 ;
        RECT 107.825 125.390 108.225 126.490 ;
        RECT 109.825 125.390 110.225 126.490 ;
        RECT 111.825 125.390 112.225 126.490 ;
        RECT 113.825 125.390 114.225 126.490 ;
        RECT 115.825 125.390 116.225 126.490 ;
        RECT 117.825 125.390 118.225 126.490 ;
        RECT 119.825 125.390 120.225 126.490 ;
        RECT 121.825 125.390 122.225 126.490 ;
        RECT 123.825 125.390 124.225 126.490 ;
        RECT 125.825 125.390 126.225 126.490 ;
        RECT 127.825 125.390 128.225 126.490 ;
        RECT 129.825 125.390 130.225 126.490 ;
        RECT 131.825 125.390 132.225 126.490 ;
        RECT 133.825 125.390 134.225 126.490 ;
        RECT 135.825 125.390 136.225 126.490 ;
        RECT 137.825 125.390 138.225 126.490 ;
        RECT 139.825 125.390 140.225 126.490 ;
        RECT 141.825 125.390 142.225 126.490 ;
        RECT 143.825 125.390 144.225 126.490 ;
        RECT 145.825 125.390 146.225 126.490 ;
        RECT 147.825 125.390 148.225 126.490 ;
        RECT 149.825 125.390 150.225 126.490 ;
        RECT 151.825 125.390 152.225 126.490 ;
        RECT 153.825 125.390 154.225 126.490 ;
        RECT 87.825 123.540 88.225 124.640 ;
        RECT 89.825 123.540 90.225 124.640 ;
        RECT 91.825 123.540 92.225 124.640 ;
        RECT 93.825 123.540 94.225 124.640 ;
        RECT 95.825 123.540 96.225 124.640 ;
        RECT 97.825 123.540 98.225 124.640 ;
        RECT 99.825 123.540 100.225 124.640 ;
        RECT 101.825 123.540 102.225 124.640 ;
        RECT 103.825 123.540 104.225 124.640 ;
        RECT 105.825 123.540 106.225 124.640 ;
        RECT 107.825 123.540 108.225 124.640 ;
        RECT 109.825 123.540 110.225 124.640 ;
        RECT 111.825 123.540 112.225 124.640 ;
        RECT 113.825 123.540 114.225 124.640 ;
        RECT 115.825 123.540 116.225 124.640 ;
        RECT 117.825 123.540 118.225 124.640 ;
        RECT 119.825 123.540 120.225 124.640 ;
        RECT 121.825 123.540 122.225 124.640 ;
        RECT 123.825 123.540 124.225 124.640 ;
        RECT 125.825 123.540 126.225 124.640 ;
        RECT 127.825 123.540 128.225 124.640 ;
        RECT 129.825 123.540 130.225 124.640 ;
        RECT 131.825 123.540 132.225 124.640 ;
        RECT 133.825 123.540 134.225 124.640 ;
        RECT 135.825 123.540 136.225 124.640 ;
        RECT 137.825 123.540 138.225 124.640 ;
        RECT 139.825 123.540 140.225 124.640 ;
        RECT 141.825 123.540 142.225 124.640 ;
        RECT 143.825 123.540 144.225 124.640 ;
        RECT 145.825 123.540 146.225 124.640 ;
        RECT 147.825 123.540 148.225 124.640 ;
        RECT 149.825 123.540 150.225 124.640 ;
        RECT 151.825 123.540 152.225 124.640 ;
        RECT 153.825 123.540 154.225 124.640 ;
        RECT 87.825 121.690 88.225 122.790 ;
        RECT 89.825 121.690 90.225 122.790 ;
        RECT 91.825 121.690 92.225 122.790 ;
        RECT 93.825 121.690 94.225 122.790 ;
        RECT 95.825 121.690 96.225 122.790 ;
        RECT 97.825 121.690 98.225 122.790 ;
        RECT 99.825 121.690 100.225 122.790 ;
        RECT 101.825 121.690 102.225 122.790 ;
        RECT 103.825 121.690 104.225 122.790 ;
        RECT 105.825 121.690 106.225 122.790 ;
        RECT 107.825 121.690 108.225 122.790 ;
        RECT 109.825 121.690 110.225 122.790 ;
        RECT 111.825 121.690 112.225 122.790 ;
        RECT 113.825 121.690 114.225 122.790 ;
        RECT 115.825 121.690 116.225 122.790 ;
        RECT 117.825 121.690 118.225 122.790 ;
        RECT 119.825 121.690 120.225 122.790 ;
        RECT 121.825 121.690 122.225 122.790 ;
        RECT 123.825 121.690 124.225 122.790 ;
        RECT 125.825 121.690 126.225 122.790 ;
        RECT 127.825 121.690 128.225 122.790 ;
        RECT 129.825 121.690 130.225 122.790 ;
        RECT 131.825 121.690 132.225 122.790 ;
        RECT 133.825 121.690 134.225 122.790 ;
        RECT 135.825 121.690 136.225 122.790 ;
        RECT 137.825 121.690 138.225 122.790 ;
        RECT 139.825 121.690 140.225 122.790 ;
        RECT 141.825 121.690 142.225 122.790 ;
        RECT 143.825 121.690 144.225 122.790 ;
        RECT 145.825 121.690 146.225 122.790 ;
        RECT 147.825 121.690 148.225 122.790 ;
        RECT 149.825 121.690 150.225 122.790 ;
        RECT 151.825 121.690 152.225 122.790 ;
        RECT 153.825 121.690 154.225 122.790 ;
        RECT 87.825 119.840 88.225 120.940 ;
        RECT 89.825 119.840 90.225 120.940 ;
        RECT 91.825 119.840 92.225 120.940 ;
        RECT 93.825 119.840 94.225 120.940 ;
        RECT 95.825 119.840 96.225 120.940 ;
        RECT 97.825 119.840 98.225 120.940 ;
        RECT 99.825 119.840 100.225 120.940 ;
        RECT 101.825 119.840 102.225 120.940 ;
        RECT 103.825 119.840 104.225 120.940 ;
        RECT 105.825 119.840 106.225 120.940 ;
        RECT 107.825 119.840 108.225 120.940 ;
        RECT 109.825 119.840 110.225 120.940 ;
        RECT 111.825 119.840 112.225 120.940 ;
        RECT 113.825 119.840 114.225 120.940 ;
        RECT 115.825 119.840 116.225 120.940 ;
        RECT 117.825 119.840 118.225 120.940 ;
        RECT 119.825 119.840 120.225 120.940 ;
        RECT 121.825 119.840 122.225 120.940 ;
        RECT 123.825 119.840 124.225 120.940 ;
        RECT 125.825 119.840 126.225 120.940 ;
        RECT 127.825 119.840 128.225 120.940 ;
        RECT 129.825 119.840 130.225 120.940 ;
        RECT 131.825 119.840 132.225 120.940 ;
        RECT 133.825 119.840 134.225 120.940 ;
        RECT 135.825 119.840 136.225 120.940 ;
        RECT 137.825 119.840 138.225 120.940 ;
        RECT 139.825 119.840 140.225 120.940 ;
        RECT 141.825 119.840 142.225 120.940 ;
        RECT 143.825 119.840 144.225 120.940 ;
        RECT 145.825 119.840 146.225 120.940 ;
        RECT 147.825 119.840 148.225 120.940 ;
        RECT 149.825 119.840 150.225 120.940 ;
        RECT 151.825 119.840 152.225 120.940 ;
        RECT 153.825 119.840 154.225 120.940 ;
        RECT 87.825 117.990 88.225 119.090 ;
        RECT 89.825 117.990 90.225 119.090 ;
        RECT 91.825 117.990 92.225 119.090 ;
        RECT 93.825 117.990 94.225 119.090 ;
        RECT 95.825 117.990 96.225 119.090 ;
        RECT 97.825 117.990 98.225 119.090 ;
        RECT 99.825 117.990 100.225 119.090 ;
        RECT 101.825 117.990 102.225 119.090 ;
        RECT 103.825 117.990 104.225 119.090 ;
        RECT 105.825 117.990 106.225 119.090 ;
        RECT 107.825 117.990 108.225 119.090 ;
        RECT 109.825 117.990 110.225 119.090 ;
        RECT 111.825 117.990 112.225 119.090 ;
        RECT 113.825 117.990 114.225 119.090 ;
        RECT 115.825 117.990 116.225 119.090 ;
        RECT 117.825 117.990 118.225 119.090 ;
        RECT 119.825 117.990 120.225 119.090 ;
        RECT 121.825 117.990 122.225 119.090 ;
        RECT 123.825 117.990 124.225 119.090 ;
        RECT 125.825 117.990 126.225 119.090 ;
        RECT 127.825 117.990 128.225 119.090 ;
        RECT 129.825 117.990 130.225 119.090 ;
        RECT 131.825 117.990 132.225 119.090 ;
        RECT 133.825 117.990 134.225 119.090 ;
        RECT 135.825 117.990 136.225 119.090 ;
        RECT 137.825 117.990 138.225 119.090 ;
        RECT 139.825 117.990 140.225 119.090 ;
        RECT 141.825 117.990 142.225 119.090 ;
        RECT 143.825 117.990 144.225 119.090 ;
        RECT 145.825 117.990 146.225 119.090 ;
        RECT 147.825 117.990 148.225 119.090 ;
        RECT 149.825 117.990 150.225 119.090 ;
        RECT 151.825 117.990 152.225 119.090 ;
        RECT 153.825 117.990 154.225 119.090 ;
        RECT 87.825 116.140 88.225 117.240 ;
        RECT 89.825 116.140 90.225 117.240 ;
        RECT 91.825 116.140 92.225 117.240 ;
        RECT 93.825 116.140 94.225 117.240 ;
        RECT 95.825 116.140 96.225 117.240 ;
        RECT 97.825 116.140 98.225 117.240 ;
        RECT 99.825 116.140 100.225 117.240 ;
        RECT 101.825 116.140 102.225 117.240 ;
        RECT 103.825 116.140 104.225 117.240 ;
        RECT 105.825 116.140 106.225 117.240 ;
        RECT 107.825 116.140 108.225 117.240 ;
        RECT 109.825 116.140 110.225 117.240 ;
        RECT 111.825 116.140 112.225 117.240 ;
        RECT 113.825 116.140 114.225 117.240 ;
        RECT 115.825 116.140 116.225 117.240 ;
        RECT 117.825 116.140 118.225 117.240 ;
        RECT 119.825 116.140 120.225 117.240 ;
        RECT 121.825 116.140 122.225 117.240 ;
        RECT 123.825 116.140 124.225 117.240 ;
        RECT 125.825 116.140 126.225 117.240 ;
        RECT 127.825 116.140 128.225 117.240 ;
        RECT 129.825 116.140 130.225 117.240 ;
        RECT 131.825 116.140 132.225 117.240 ;
        RECT 133.825 116.140 134.225 117.240 ;
        RECT 135.825 116.140 136.225 117.240 ;
        RECT 137.825 116.140 138.225 117.240 ;
        RECT 139.825 116.140 140.225 117.240 ;
        RECT 141.825 116.140 142.225 117.240 ;
        RECT 143.825 116.140 144.225 117.240 ;
        RECT 145.825 116.140 146.225 117.240 ;
        RECT 147.825 116.140 148.225 117.240 ;
        RECT 149.825 116.140 150.225 117.240 ;
        RECT 151.825 116.140 152.225 117.240 ;
        RECT 153.825 116.140 154.225 117.240 ;
        RECT 87.825 114.290 88.225 115.390 ;
        RECT 89.825 114.290 90.225 115.390 ;
        RECT 91.825 114.290 92.225 115.390 ;
        RECT 93.825 114.290 94.225 115.390 ;
        RECT 95.825 114.290 96.225 115.390 ;
        RECT 97.825 114.290 98.225 115.390 ;
        RECT 99.825 114.290 100.225 115.390 ;
        RECT 101.825 114.290 102.225 115.390 ;
        RECT 103.825 114.290 104.225 115.390 ;
        RECT 105.825 114.290 106.225 115.390 ;
        RECT 107.825 114.290 108.225 115.390 ;
        RECT 109.825 114.290 110.225 115.390 ;
        RECT 111.825 114.290 112.225 115.390 ;
        RECT 113.825 114.290 114.225 115.390 ;
        RECT 115.825 114.290 116.225 115.390 ;
        RECT 117.825 114.290 118.225 115.390 ;
        RECT 119.825 114.290 120.225 115.390 ;
        RECT 121.825 114.290 122.225 115.390 ;
        RECT 123.825 114.290 124.225 115.390 ;
        RECT 125.825 114.290 126.225 115.390 ;
        RECT 127.825 114.290 128.225 115.390 ;
        RECT 129.825 114.290 130.225 115.390 ;
        RECT 131.825 114.290 132.225 115.390 ;
        RECT 133.825 114.290 134.225 115.390 ;
        RECT 135.825 114.290 136.225 115.390 ;
        RECT 137.825 114.290 138.225 115.390 ;
        RECT 139.825 114.290 140.225 115.390 ;
        RECT 141.825 114.290 142.225 115.390 ;
        RECT 143.825 114.290 144.225 115.390 ;
        RECT 145.825 114.290 146.225 115.390 ;
        RECT 147.825 114.290 148.225 115.390 ;
        RECT 149.825 114.290 150.225 115.390 ;
        RECT 151.825 114.290 152.225 115.390 ;
        RECT 153.825 114.290 154.225 115.390 ;
        RECT 87.825 112.440 88.225 113.540 ;
        RECT 89.825 112.440 90.225 113.540 ;
        RECT 91.825 112.440 92.225 113.540 ;
        RECT 93.825 112.440 94.225 113.540 ;
        RECT 95.825 112.440 96.225 113.540 ;
        RECT 97.825 112.440 98.225 113.540 ;
        RECT 99.825 112.440 100.225 113.540 ;
        RECT 101.825 112.440 102.225 113.540 ;
        RECT 103.825 112.440 104.225 113.540 ;
        RECT 105.825 112.440 106.225 113.540 ;
        RECT 107.825 112.440 108.225 113.540 ;
        RECT 109.825 112.440 110.225 113.540 ;
        RECT 111.825 112.440 112.225 113.540 ;
        RECT 113.825 112.440 114.225 113.540 ;
        RECT 115.825 112.440 116.225 113.540 ;
        RECT 117.825 112.440 118.225 113.540 ;
        RECT 119.825 112.440 120.225 113.540 ;
        RECT 121.825 112.440 122.225 113.540 ;
        RECT 123.825 112.440 124.225 113.540 ;
        RECT 125.825 112.440 126.225 113.540 ;
        RECT 127.825 112.440 128.225 113.540 ;
        RECT 129.825 112.440 130.225 113.540 ;
        RECT 131.825 112.440 132.225 113.540 ;
        RECT 133.825 112.440 134.225 113.540 ;
        RECT 135.825 112.440 136.225 113.540 ;
        RECT 137.825 112.440 138.225 113.540 ;
        RECT 139.825 112.440 140.225 113.540 ;
        RECT 141.825 112.440 142.225 113.540 ;
        RECT 143.825 112.440 144.225 113.540 ;
        RECT 145.825 112.440 146.225 113.540 ;
        RECT 147.825 112.440 148.225 113.540 ;
        RECT 149.825 112.440 150.225 113.540 ;
        RECT 151.825 112.440 152.225 113.540 ;
        RECT 153.825 112.440 154.225 113.540 ;
        RECT 87.825 110.590 88.225 111.690 ;
        RECT 89.825 110.590 90.225 111.690 ;
        RECT 91.825 110.590 92.225 111.690 ;
        RECT 93.825 110.590 94.225 111.690 ;
        RECT 95.825 110.590 96.225 111.690 ;
        RECT 97.825 110.590 98.225 111.690 ;
        RECT 99.825 110.590 100.225 111.690 ;
        RECT 101.825 110.590 102.225 111.690 ;
        RECT 103.825 110.590 104.225 111.690 ;
        RECT 105.825 110.590 106.225 111.690 ;
        RECT 107.825 110.590 108.225 111.690 ;
        RECT 109.825 110.590 110.225 111.690 ;
        RECT 111.825 110.590 112.225 111.690 ;
        RECT 113.825 110.590 114.225 111.690 ;
        RECT 115.825 110.590 116.225 111.690 ;
        RECT 117.825 110.590 118.225 111.690 ;
        RECT 119.825 110.590 120.225 111.690 ;
        RECT 121.825 110.590 122.225 111.690 ;
        RECT 123.825 110.590 124.225 111.690 ;
        RECT 125.825 110.590 126.225 111.690 ;
        RECT 127.825 110.590 128.225 111.690 ;
        RECT 129.825 110.590 130.225 111.690 ;
        RECT 131.825 110.590 132.225 111.690 ;
        RECT 133.825 110.590 134.225 111.690 ;
        RECT 135.825 110.590 136.225 111.690 ;
        RECT 137.825 110.590 138.225 111.690 ;
        RECT 139.825 110.590 140.225 111.690 ;
        RECT 141.825 110.590 142.225 111.690 ;
        RECT 143.825 110.590 144.225 111.690 ;
        RECT 145.825 110.590 146.225 111.690 ;
        RECT 147.825 110.590 148.225 111.690 ;
        RECT 149.825 110.590 150.225 111.690 ;
        RECT 151.825 110.590 152.225 111.690 ;
        RECT 153.825 110.590 154.225 111.690 ;
        RECT 87.825 108.740 88.225 109.840 ;
        RECT 89.825 108.740 90.225 109.840 ;
        RECT 91.825 108.740 92.225 109.840 ;
        RECT 93.825 108.740 94.225 109.840 ;
        RECT 95.825 108.740 96.225 109.840 ;
        RECT 97.825 108.740 98.225 109.840 ;
        RECT 99.825 108.740 100.225 109.840 ;
        RECT 101.825 108.740 102.225 109.840 ;
        RECT 103.825 108.740 104.225 109.840 ;
        RECT 105.825 108.740 106.225 109.840 ;
        RECT 107.825 108.740 108.225 109.840 ;
        RECT 109.825 108.740 110.225 109.840 ;
        RECT 111.825 108.740 112.225 109.840 ;
        RECT 113.825 108.740 114.225 109.840 ;
        RECT 115.825 108.740 116.225 109.840 ;
        RECT 117.825 108.740 118.225 109.840 ;
        RECT 119.825 108.740 120.225 109.840 ;
        RECT 121.825 108.740 122.225 109.840 ;
        RECT 123.825 108.740 124.225 109.840 ;
        RECT 125.825 108.740 126.225 109.840 ;
        RECT 127.825 108.740 128.225 109.840 ;
        RECT 129.825 108.740 130.225 109.840 ;
        RECT 131.825 108.740 132.225 109.840 ;
        RECT 133.825 108.740 134.225 109.840 ;
        RECT 135.825 108.740 136.225 109.840 ;
        RECT 137.825 108.740 138.225 109.840 ;
        RECT 139.825 108.740 140.225 109.840 ;
        RECT 141.825 108.740 142.225 109.840 ;
        RECT 143.825 108.740 144.225 109.840 ;
        RECT 145.825 108.740 146.225 109.840 ;
        RECT 147.825 108.740 148.225 109.840 ;
        RECT 149.825 108.740 150.225 109.840 ;
        RECT 151.825 108.740 152.225 109.840 ;
        RECT 153.825 108.740 154.225 109.840 ;
        RECT 87.825 106.890 88.225 107.990 ;
        RECT 89.825 106.890 90.225 107.990 ;
        RECT 91.825 106.890 92.225 107.990 ;
        RECT 93.825 106.890 94.225 107.990 ;
        RECT 95.825 106.890 96.225 107.990 ;
        RECT 97.825 106.890 98.225 107.990 ;
        RECT 99.825 106.890 100.225 107.990 ;
        RECT 101.825 106.890 102.225 107.990 ;
        RECT 103.825 106.890 104.225 107.990 ;
        RECT 105.825 106.890 106.225 107.990 ;
        RECT 107.825 106.890 108.225 107.990 ;
        RECT 109.825 106.890 110.225 107.990 ;
        RECT 111.825 106.890 112.225 107.990 ;
        RECT 113.825 106.890 114.225 107.990 ;
        RECT 115.825 106.890 116.225 107.990 ;
        RECT 117.825 106.890 118.225 107.990 ;
        RECT 119.825 106.890 120.225 107.990 ;
        RECT 121.825 106.890 122.225 107.990 ;
        RECT 123.825 106.890 124.225 107.990 ;
        RECT 125.825 106.890 126.225 107.990 ;
        RECT 127.825 106.890 128.225 107.990 ;
        RECT 129.825 106.890 130.225 107.990 ;
        RECT 131.825 106.890 132.225 107.990 ;
        RECT 133.825 106.890 134.225 107.990 ;
        RECT 135.825 106.890 136.225 107.990 ;
        RECT 137.825 106.890 138.225 107.990 ;
        RECT 139.825 106.890 140.225 107.990 ;
        RECT 141.825 106.890 142.225 107.990 ;
        RECT 143.825 106.890 144.225 107.990 ;
        RECT 145.825 106.890 146.225 107.990 ;
        RECT 147.825 106.890 148.225 107.990 ;
        RECT 149.825 106.890 150.225 107.990 ;
        RECT 151.825 106.890 152.225 107.990 ;
        RECT 153.825 106.890 154.225 107.990 ;
        RECT 87.825 105.040 88.225 106.140 ;
        RECT 89.825 105.040 90.225 106.140 ;
        RECT 91.825 105.040 92.225 106.140 ;
        RECT 93.825 105.040 94.225 106.140 ;
        RECT 95.825 105.040 96.225 106.140 ;
        RECT 97.825 105.040 98.225 106.140 ;
        RECT 99.825 105.040 100.225 106.140 ;
        RECT 101.825 105.040 102.225 106.140 ;
        RECT 103.825 105.040 104.225 106.140 ;
        RECT 105.825 105.040 106.225 106.140 ;
        RECT 107.825 105.040 108.225 106.140 ;
        RECT 109.825 105.040 110.225 106.140 ;
        RECT 111.825 105.040 112.225 106.140 ;
        RECT 113.825 105.040 114.225 106.140 ;
        RECT 115.825 105.040 116.225 106.140 ;
        RECT 117.825 105.040 118.225 106.140 ;
        RECT 119.825 105.040 120.225 106.140 ;
        RECT 121.825 105.040 122.225 106.140 ;
        RECT 123.825 105.040 124.225 106.140 ;
        RECT 125.825 105.040 126.225 106.140 ;
        RECT 127.825 105.040 128.225 106.140 ;
        RECT 129.825 105.040 130.225 106.140 ;
        RECT 131.825 105.040 132.225 106.140 ;
        RECT 133.825 105.040 134.225 106.140 ;
        RECT 135.825 105.040 136.225 106.140 ;
        RECT 137.825 105.040 138.225 106.140 ;
        RECT 139.825 105.040 140.225 106.140 ;
        RECT 141.825 105.040 142.225 106.140 ;
        RECT 143.825 105.040 144.225 106.140 ;
        RECT 145.825 105.040 146.225 106.140 ;
        RECT 147.825 105.040 148.225 106.140 ;
        RECT 149.825 105.040 150.225 106.140 ;
        RECT 151.825 105.040 152.225 106.140 ;
        RECT 153.825 105.040 154.225 106.140 ;
        RECT 87.825 103.190 88.225 104.290 ;
        RECT 89.825 103.190 90.225 104.290 ;
        RECT 91.825 103.190 92.225 104.290 ;
        RECT 93.825 103.190 94.225 104.290 ;
        RECT 95.825 103.190 96.225 104.290 ;
        RECT 97.825 103.190 98.225 104.290 ;
        RECT 99.825 103.190 100.225 104.290 ;
        RECT 101.825 103.190 102.225 104.290 ;
        RECT 103.825 103.190 104.225 104.290 ;
        RECT 105.825 103.190 106.225 104.290 ;
        RECT 107.825 103.190 108.225 104.290 ;
        RECT 109.825 103.190 110.225 104.290 ;
        RECT 111.825 103.190 112.225 104.290 ;
        RECT 113.825 103.190 114.225 104.290 ;
        RECT 115.825 103.190 116.225 104.290 ;
        RECT 117.825 103.190 118.225 104.290 ;
        RECT 119.825 103.190 120.225 104.290 ;
        RECT 121.825 103.190 122.225 104.290 ;
        RECT 123.825 103.190 124.225 104.290 ;
        RECT 125.825 103.190 126.225 104.290 ;
        RECT 127.825 103.190 128.225 104.290 ;
        RECT 129.825 103.190 130.225 104.290 ;
        RECT 131.825 103.190 132.225 104.290 ;
        RECT 133.825 103.190 134.225 104.290 ;
        RECT 135.825 103.190 136.225 104.290 ;
        RECT 137.825 103.190 138.225 104.290 ;
        RECT 139.825 103.190 140.225 104.290 ;
        RECT 141.825 103.190 142.225 104.290 ;
        RECT 143.825 103.190 144.225 104.290 ;
        RECT 145.825 103.190 146.225 104.290 ;
        RECT 147.825 103.190 148.225 104.290 ;
        RECT 149.825 103.190 150.225 104.290 ;
        RECT 151.825 103.190 152.225 104.290 ;
        RECT 153.825 103.190 154.225 104.290 ;
        RECT 87.825 101.340 88.225 102.440 ;
        RECT 89.825 101.340 90.225 102.440 ;
        RECT 91.825 101.340 92.225 102.440 ;
        RECT 93.825 101.340 94.225 102.440 ;
        RECT 95.825 101.340 96.225 102.440 ;
        RECT 97.825 101.340 98.225 102.440 ;
        RECT 99.825 101.340 100.225 102.440 ;
        RECT 101.825 101.340 102.225 102.440 ;
        RECT 103.825 101.340 104.225 102.440 ;
        RECT 105.825 101.340 106.225 102.440 ;
        RECT 107.825 101.340 108.225 102.440 ;
        RECT 109.825 101.340 110.225 102.440 ;
        RECT 111.825 101.340 112.225 102.440 ;
        RECT 113.825 101.340 114.225 102.440 ;
        RECT 115.825 101.340 116.225 102.440 ;
        RECT 117.825 101.340 118.225 102.440 ;
        RECT 119.825 101.340 120.225 102.440 ;
        RECT 121.825 101.340 122.225 102.440 ;
        RECT 123.825 101.340 124.225 102.440 ;
        RECT 125.825 101.340 126.225 102.440 ;
        RECT 127.825 101.340 128.225 102.440 ;
        RECT 129.825 101.340 130.225 102.440 ;
        RECT 131.825 101.340 132.225 102.440 ;
        RECT 133.825 101.340 134.225 102.440 ;
        RECT 135.825 101.340 136.225 102.440 ;
        RECT 137.825 101.340 138.225 102.440 ;
        RECT 139.825 101.340 140.225 102.440 ;
        RECT 141.825 101.340 142.225 102.440 ;
        RECT 143.825 101.340 144.225 102.440 ;
        RECT 145.825 101.340 146.225 102.440 ;
        RECT 147.825 101.340 148.225 102.440 ;
        RECT 149.825 101.340 150.225 102.440 ;
        RECT 151.825 101.340 152.225 102.440 ;
        RECT 153.825 101.340 154.225 102.440 ;
        RECT 87.825 99.490 88.225 100.590 ;
        RECT 89.825 99.490 90.225 100.590 ;
        RECT 91.825 99.490 92.225 100.590 ;
        RECT 93.825 99.490 94.225 100.590 ;
        RECT 95.825 99.490 96.225 100.590 ;
        RECT 97.825 99.490 98.225 100.590 ;
        RECT 99.825 99.490 100.225 100.590 ;
        RECT 101.825 99.490 102.225 100.590 ;
        RECT 103.825 99.490 104.225 100.590 ;
        RECT 105.825 99.490 106.225 100.590 ;
        RECT 107.825 99.490 108.225 100.590 ;
        RECT 109.825 99.490 110.225 100.590 ;
        RECT 111.825 99.490 112.225 100.590 ;
        RECT 113.825 99.490 114.225 100.590 ;
        RECT 115.825 99.490 116.225 100.590 ;
        RECT 117.825 99.490 118.225 100.590 ;
        RECT 119.825 99.490 120.225 100.590 ;
        RECT 121.825 99.490 122.225 100.590 ;
        RECT 123.825 99.490 124.225 100.590 ;
        RECT 125.825 99.490 126.225 100.590 ;
        RECT 127.825 99.490 128.225 100.590 ;
        RECT 129.825 99.490 130.225 100.590 ;
        RECT 131.825 99.490 132.225 100.590 ;
        RECT 133.825 99.490 134.225 100.590 ;
        RECT 135.825 99.490 136.225 100.590 ;
        RECT 137.825 99.490 138.225 100.590 ;
        RECT 139.825 99.490 140.225 100.590 ;
        RECT 141.825 99.490 142.225 100.590 ;
        RECT 143.825 99.490 144.225 100.590 ;
        RECT 145.825 99.490 146.225 100.590 ;
        RECT 147.825 99.490 148.225 100.590 ;
        RECT 149.825 99.490 150.225 100.590 ;
        RECT 151.825 99.490 152.225 100.590 ;
        RECT 153.825 99.490 154.225 100.590 ;
        RECT 87.825 97.640 88.225 98.740 ;
        RECT 89.825 97.640 90.225 98.740 ;
        RECT 91.825 97.640 92.225 98.740 ;
        RECT 93.825 97.640 94.225 98.740 ;
        RECT 95.825 97.640 96.225 98.740 ;
        RECT 97.825 97.640 98.225 98.740 ;
        RECT 99.825 97.640 100.225 98.740 ;
        RECT 101.825 97.640 102.225 98.740 ;
        RECT 103.825 97.640 104.225 98.740 ;
        RECT 105.825 97.640 106.225 98.740 ;
        RECT 107.825 97.640 108.225 98.740 ;
        RECT 109.825 97.640 110.225 98.740 ;
        RECT 111.825 97.640 112.225 98.740 ;
        RECT 113.825 97.640 114.225 98.740 ;
        RECT 115.825 97.640 116.225 98.740 ;
        RECT 117.825 97.640 118.225 98.740 ;
        RECT 119.825 97.640 120.225 98.740 ;
        RECT 121.825 97.640 122.225 98.740 ;
        RECT 123.825 97.640 124.225 98.740 ;
        RECT 125.825 97.640 126.225 98.740 ;
        RECT 127.825 97.640 128.225 98.740 ;
        RECT 129.825 97.640 130.225 98.740 ;
        RECT 131.825 97.640 132.225 98.740 ;
        RECT 133.825 97.640 134.225 98.740 ;
        RECT 135.825 97.640 136.225 98.740 ;
        RECT 137.825 97.640 138.225 98.740 ;
        RECT 139.825 97.640 140.225 98.740 ;
        RECT 141.825 97.640 142.225 98.740 ;
        RECT 143.825 97.640 144.225 98.740 ;
        RECT 145.825 97.640 146.225 98.740 ;
        RECT 147.825 97.640 148.225 98.740 ;
        RECT 149.825 97.640 150.225 98.740 ;
        RECT 151.825 97.640 152.225 98.740 ;
        RECT 153.825 97.640 154.225 98.740 ;
        RECT 87.825 95.790 88.225 96.890 ;
        RECT 89.825 95.790 90.225 96.890 ;
        RECT 91.825 95.790 92.225 96.890 ;
        RECT 93.825 95.790 94.225 96.890 ;
        RECT 95.825 95.790 96.225 96.890 ;
        RECT 97.825 95.790 98.225 96.890 ;
        RECT 99.825 95.790 100.225 96.890 ;
        RECT 101.825 95.790 102.225 96.890 ;
        RECT 103.825 95.790 104.225 96.890 ;
        RECT 105.825 95.790 106.225 96.890 ;
        RECT 107.825 95.790 108.225 96.890 ;
        RECT 109.825 95.790 110.225 96.890 ;
        RECT 111.825 95.790 112.225 96.890 ;
        RECT 113.825 95.790 114.225 96.890 ;
        RECT 115.825 95.790 116.225 96.890 ;
        RECT 117.825 95.790 118.225 96.890 ;
        RECT 119.825 95.790 120.225 96.890 ;
        RECT 121.825 95.790 122.225 96.890 ;
        RECT 123.825 95.790 124.225 96.890 ;
        RECT 125.825 95.790 126.225 96.890 ;
        RECT 127.825 95.790 128.225 96.890 ;
        RECT 129.825 95.790 130.225 96.890 ;
        RECT 131.825 95.790 132.225 96.890 ;
        RECT 133.825 95.790 134.225 96.890 ;
        RECT 135.825 95.790 136.225 96.890 ;
        RECT 137.825 95.790 138.225 96.890 ;
        RECT 139.825 95.790 140.225 96.890 ;
        RECT 141.825 95.790 142.225 96.890 ;
        RECT 143.825 95.790 144.225 96.890 ;
        RECT 145.825 95.790 146.225 96.890 ;
        RECT 147.825 95.790 148.225 96.890 ;
        RECT 149.825 95.790 150.225 96.890 ;
        RECT 151.825 95.790 152.225 96.890 ;
        RECT 153.825 95.790 154.225 96.890 ;
        RECT 87.825 93.940 88.225 95.040 ;
        RECT 89.825 93.940 90.225 95.040 ;
        RECT 91.825 93.940 92.225 95.040 ;
        RECT 93.825 93.940 94.225 95.040 ;
        RECT 95.825 93.940 96.225 95.040 ;
        RECT 97.825 93.940 98.225 95.040 ;
        RECT 99.825 93.940 100.225 95.040 ;
        RECT 101.825 93.940 102.225 95.040 ;
        RECT 103.825 93.940 104.225 95.040 ;
        RECT 105.825 93.940 106.225 95.040 ;
        RECT 107.825 93.940 108.225 95.040 ;
        RECT 109.825 93.940 110.225 95.040 ;
        RECT 111.825 93.940 112.225 95.040 ;
        RECT 113.825 93.940 114.225 95.040 ;
        RECT 115.825 93.940 116.225 95.040 ;
        RECT 117.825 93.940 118.225 95.040 ;
        RECT 119.825 93.940 120.225 95.040 ;
        RECT 121.825 93.940 122.225 95.040 ;
        RECT 123.825 93.940 124.225 95.040 ;
        RECT 125.825 93.940 126.225 95.040 ;
        RECT 127.825 93.940 128.225 95.040 ;
        RECT 129.825 93.940 130.225 95.040 ;
        RECT 131.825 93.940 132.225 95.040 ;
        RECT 133.825 93.940 134.225 95.040 ;
        RECT 135.825 93.940 136.225 95.040 ;
        RECT 137.825 93.940 138.225 95.040 ;
        RECT 139.825 93.940 140.225 95.040 ;
        RECT 141.825 93.940 142.225 95.040 ;
        RECT 143.825 93.940 144.225 95.040 ;
        RECT 145.825 93.940 146.225 95.040 ;
        RECT 147.825 93.940 148.225 95.040 ;
        RECT 149.825 93.940 150.225 95.040 ;
        RECT 151.825 93.940 152.225 95.040 ;
        RECT 153.825 93.940 154.225 95.040 ;
        RECT 87.825 92.090 88.225 93.190 ;
        RECT 89.825 92.090 90.225 93.190 ;
        RECT 91.825 92.090 92.225 93.190 ;
        RECT 93.825 92.090 94.225 93.190 ;
        RECT 95.825 92.090 96.225 93.190 ;
        RECT 97.825 92.090 98.225 93.190 ;
        RECT 99.825 92.090 100.225 93.190 ;
        RECT 101.825 92.090 102.225 93.190 ;
        RECT 103.825 92.090 104.225 93.190 ;
        RECT 105.825 92.090 106.225 93.190 ;
        RECT 107.825 92.090 108.225 93.190 ;
        RECT 109.825 92.090 110.225 93.190 ;
        RECT 111.825 92.090 112.225 93.190 ;
        RECT 113.825 92.090 114.225 93.190 ;
        RECT 115.825 92.090 116.225 93.190 ;
        RECT 117.825 92.090 118.225 93.190 ;
        RECT 119.825 92.090 120.225 93.190 ;
        RECT 121.825 92.090 122.225 93.190 ;
        RECT 123.825 92.090 124.225 93.190 ;
        RECT 125.825 92.090 126.225 93.190 ;
        RECT 127.825 92.090 128.225 93.190 ;
        RECT 129.825 92.090 130.225 93.190 ;
        RECT 131.825 92.090 132.225 93.190 ;
        RECT 133.825 92.090 134.225 93.190 ;
        RECT 135.825 92.090 136.225 93.190 ;
        RECT 137.825 92.090 138.225 93.190 ;
        RECT 139.825 92.090 140.225 93.190 ;
        RECT 141.825 92.090 142.225 93.190 ;
        RECT 143.825 92.090 144.225 93.190 ;
        RECT 145.825 92.090 146.225 93.190 ;
        RECT 147.825 92.090 148.225 93.190 ;
        RECT 149.825 92.090 150.225 93.190 ;
        RECT 151.825 92.090 152.225 93.190 ;
        RECT 153.825 92.090 154.225 93.190 ;
        RECT 87.825 90.240 88.225 91.340 ;
        RECT 89.825 90.240 90.225 91.340 ;
        RECT 91.825 90.240 92.225 91.340 ;
        RECT 93.825 90.240 94.225 91.340 ;
        RECT 95.825 90.240 96.225 91.340 ;
        RECT 97.825 90.240 98.225 91.340 ;
        RECT 99.825 90.240 100.225 91.340 ;
        RECT 101.825 90.240 102.225 91.340 ;
        RECT 103.825 90.240 104.225 91.340 ;
        RECT 105.825 90.240 106.225 91.340 ;
        RECT 107.825 90.240 108.225 91.340 ;
        RECT 109.825 90.240 110.225 91.340 ;
        RECT 111.825 90.240 112.225 91.340 ;
        RECT 113.825 90.240 114.225 91.340 ;
        RECT 115.825 90.240 116.225 91.340 ;
        RECT 117.825 90.240 118.225 91.340 ;
        RECT 119.825 90.240 120.225 91.340 ;
        RECT 121.825 90.240 122.225 91.340 ;
        RECT 123.825 90.240 124.225 91.340 ;
        RECT 125.825 90.240 126.225 91.340 ;
        RECT 127.825 90.240 128.225 91.340 ;
        RECT 129.825 90.240 130.225 91.340 ;
        RECT 131.825 90.240 132.225 91.340 ;
        RECT 133.825 90.240 134.225 91.340 ;
        RECT 135.825 90.240 136.225 91.340 ;
        RECT 137.825 90.240 138.225 91.340 ;
        RECT 139.825 90.240 140.225 91.340 ;
        RECT 141.825 90.240 142.225 91.340 ;
        RECT 143.825 90.240 144.225 91.340 ;
        RECT 145.825 90.240 146.225 91.340 ;
        RECT 147.825 90.240 148.225 91.340 ;
        RECT 149.825 90.240 150.225 91.340 ;
        RECT 151.825 90.240 152.225 91.340 ;
        RECT 153.825 90.240 154.225 91.340 ;
        RECT 87.825 88.390 88.225 89.490 ;
        RECT 89.825 88.390 90.225 89.490 ;
        RECT 91.825 88.390 92.225 89.490 ;
        RECT 93.825 88.390 94.225 89.490 ;
        RECT 95.825 88.390 96.225 89.490 ;
        RECT 97.825 88.390 98.225 89.490 ;
        RECT 99.825 88.390 100.225 89.490 ;
        RECT 101.825 88.390 102.225 89.490 ;
        RECT 103.825 88.390 104.225 89.490 ;
        RECT 105.825 88.390 106.225 89.490 ;
        RECT 107.825 88.390 108.225 89.490 ;
        RECT 109.825 88.390 110.225 89.490 ;
        RECT 111.825 88.390 112.225 89.490 ;
        RECT 113.825 88.390 114.225 89.490 ;
        RECT 115.825 88.390 116.225 89.490 ;
        RECT 117.825 88.390 118.225 89.490 ;
        RECT 119.825 88.390 120.225 89.490 ;
        RECT 121.825 88.390 122.225 89.490 ;
        RECT 123.825 88.390 124.225 89.490 ;
        RECT 125.825 88.390 126.225 89.490 ;
        RECT 127.825 88.390 128.225 89.490 ;
        RECT 129.825 88.390 130.225 89.490 ;
        RECT 131.825 88.390 132.225 89.490 ;
        RECT 133.825 88.390 134.225 89.490 ;
        RECT 135.825 88.390 136.225 89.490 ;
        RECT 137.825 88.390 138.225 89.490 ;
        RECT 139.825 88.390 140.225 89.490 ;
        RECT 141.825 88.390 142.225 89.490 ;
        RECT 143.825 88.390 144.225 89.490 ;
        RECT 145.825 88.390 146.225 89.490 ;
        RECT 147.825 88.390 148.225 89.490 ;
        RECT 149.825 88.390 150.225 89.490 ;
        RECT 151.825 88.390 152.225 89.490 ;
        RECT 153.825 88.390 154.225 89.490 ;
        RECT 87.825 86.540 88.225 87.640 ;
        RECT 89.825 86.540 90.225 87.640 ;
        RECT 91.825 86.540 92.225 87.640 ;
        RECT 93.825 86.540 94.225 87.640 ;
        RECT 95.825 86.540 96.225 87.640 ;
        RECT 97.825 86.540 98.225 87.640 ;
        RECT 99.825 86.540 100.225 87.640 ;
        RECT 101.825 86.540 102.225 87.640 ;
        RECT 103.825 86.540 104.225 87.640 ;
        RECT 105.825 86.540 106.225 87.640 ;
        RECT 107.825 86.540 108.225 87.640 ;
        RECT 109.825 86.540 110.225 87.640 ;
        RECT 111.825 86.540 112.225 87.640 ;
        RECT 113.825 86.540 114.225 87.640 ;
        RECT 115.825 86.540 116.225 87.640 ;
        RECT 117.825 86.540 118.225 87.640 ;
        RECT 119.825 86.540 120.225 87.640 ;
        RECT 121.825 86.540 122.225 87.640 ;
        RECT 123.825 86.540 124.225 87.640 ;
        RECT 125.825 86.540 126.225 87.640 ;
        RECT 127.825 86.540 128.225 87.640 ;
        RECT 129.825 86.540 130.225 87.640 ;
        RECT 131.825 86.540 132.225 87.640 ;
        RECT 133.825 86.540 134.225 87.640 ;
        RECT 135.825 86.540 136.225 87.640 ;
        RECT 137.825 86.540 138.225 87.640 ;
        RECT 139.825 86.540 140.225 87.640 ;
        RECT 141.825 86.540 142.225 87.640 ;
        RECT 143.825 86.540 144.225 87.640 ;
        RECT 145.825 86.540 146.225 87.640 ;
        RECT 147.825 86.540 148.225 87.640 ;
        RECT 149.825 86.540 150.225 87.640 ;
        RECT 151.825 86.540 152.225 87.640 ;
        RECT 153.825 86.540 154.225 87.640 ;
        RECT 87.825 84.690 88.225 85.790 ;
        RECT 89.825 84.690 90.225 85.790 ;
        RECT 91.825 84.690 92.225 85.790 ;
        RECT 93.825 84.690 94.225 85.790 ;
        RECT 95.825 84.690 96.225 85.790 ;
        RECT 97.825 84.690 98.225 85.790 ;
        RECT 99.825 84.690 100.225 85.790 ;
        RECT 101.825 84.690 102.225 85.790 ;
        RECT 103.825 84.690 104.225 85.790 ;
        RECT 105.825 84.690 106.225 85.790 ;
        RECT 107.825 84.690 108.225 85.790 ;
        RECT 109.825 84.690 110.225 85.790 ;
        RECT 111.825 84.690 112.225 85.790 ;
        RECT 113.825 84.690 114.225 85.790 ;
        RECT 115.825 84.690 116.225 85.790 ;
        RECT 117.825 84.690 118.225 85.790 ;
        RECT 119.825 84.690 120.225 85.790 ;
        RECT 121.825 84.690 122.225 85.790 ;
        RECT 123.825 84.690 124.225 85.790 ;
        RECT 125.825 84.690 126.225 85.790 ;
        RECT 127.825 84.690 128.225 85.790 ;
        RECT 129.825 84.690 130.225 85.790 ;
        RECT 131.825 84.690 132.225 85.790 ;
        RECT 133.825 84.690 134.225 85.790 ;
        RECT 135.825 84.690 136.225 85.790 ;
        RECT 137.825 84.690 138.225 85.790 ;
        RECT 139.825 84.690 140.225 85.790 ;
        RECT 141.825 84.690 142.225 85.790 ;
        RECT 143.825 84.690 144.225 85.790 ;
        RECT 145.825 84.690 146.225 85.790 ;
        RECT 147.825 84.690 148.225 85.790 ;
        RECT 149.825 84.690 150.225 85.790 ;
        RECT 151.825 84.690 152.225 85.790 ;
        RECT 153.825 84.690 154.225 85.790 ;
        RECT 87.825 82.840 88.225 83.940 ;
        RECT 89.825 82.840 90.225 83.940 ;
        RECT 91.825 82.840 92.225 83.940 ;
        RECT 93.825 82.840 94.225 83.940 ;
        RECT 95.825 82.840 96.225 83.940 ;
        RECT 97.825 82.840 98.225 83.940 ;
        RECT 99.825 82.840 100.225 83.940 ;
        RECT 101.825 82.840 102.225 83.940 ;
        RECT 103.825 82.840 104.225 83.940 ;
        RECT 105.825 82.840 106.225 83.940 ;
        RECT 107.825 82.840 108.225 83.940 ;
        RECT 109.825 82.840 110.225 83.940 ;
        RECT 111.825 82.840 112.225 83.940 ;
        RECT 113.825 82.840 114.225 83.940 ;
        RECT 115.825 82.840 116.225 83.940 ;
        RECT 117.825 82.840 118.225 83.940 ;
        RECT 119.825 82.840 120.225 83.940 ;
        RECT 121.825 82.840 122.225 83.940 ;
        RECT 123.825 82.840 124.225 83.940 ;
        RECT 125.825 82.840 126.225 83.940 ;
        RECT 127.825 82.840 128.225 83.940 ;
        RECT 129.825 82.840 130.225 83.940 ;
        RECT 131.825 82.840 132.225 83.940 ;
        RECT 133.825 82.840 134.225 83.940 ;
        RECT 135.825 82.840 136.225 83.940 ;
        RECT 137.825 82.840 138.225 83.940 ;
        RECT 139.825 82.840 140.225 83.940 ;
        RECT 141.825 82.840 142.225 83.940 ;
        RECT 143.825 82.840 144.225 83.940 ;
        RECT 145.825 82.840 146.225 83.940 ;
        RECT 147.825 82.840 148.225 83.940 ;
        RECT 149.825 82.840 150.225 83.940 ;
        RECT 151.825 82.840 152.225 83.940 ;
        RECT 153.825 82.840 154.225 83.940 ;
        RECT 87.825 80.990 88.225 82.090 ;
        RECT 89.825 80.990 90.225 82.090 ;
        RECT 91.825 80.990 92.225 82.090 ;
        RECT 93.825 80.990 94.225 82.090 ;
        RECT 95.825 80.990 96.225 82.090 ;
        RECT 97.825 80.990 98.225 82.090 ;
        RECT 99.825 80.990 100.225 82.090 ;
        RECT 101.825 80.990 102.225 82.090 ;
        RECT 103.825 80.990 104.225 82.090 ;
        RECT 105.825 80.990 106.225 82.090 ;
        RECT 107.825 80.990 108.225 82.090 ;
        RECT 109.825 80.990 110.225 82.090 ;
        RECT 111.825 80.990 112.225 82.090 ;
        RECT 113.825 80.990 114.225 82.090 ;
        RECT 115.825 80.990 116.225 82.090 ;
        RECT 117.825 80.990 118.225 82.090 ;
        RECT 119.825 80.990 120.225 82.090 ;
        RECT 121.825 80.990 122.225 82.090 ;
        RECT 123.825 80.990 124.225 82.090 ;
        RECT 125.825 80.990 126.225 82.090 ;
        RECT 127.825 80.990 128.225 82.090 ;
        RECT 129.825 80.990 130.225 82.090 ;
        RECT 131.825 80.990 132.225 82.090 ;
        RECT 133.825 80.990 134.225 82.090 ;
        RECT 135.825 80.990 136.225 82.090 ;
        RECT 137.825 80.990 138.225 82.090 ;
        RECT 139.825 80.990 140.225 82.090 ;
        RECT 141.825 80.990 142.225 82.090 ;
        RECT 143.825 80.990 144.225 82.090 ;
        RECT 145.825 80.990 146.225 82.090 ;
        RECT 147.825 80.990 148.225 82.090 ;
        RECT 149.825 80.990 150.225 82.090 ;
        RECT 151.825 80.990 152.225 82.090 ;
        RECT 153.825 80.990 154.225 82.090 ;
        RECT 87.825 79.140 88.225 80.240 ;
        RECT 89.825 79.140 90.225 80.240 ;
        RECT 91.825 79.140 92.225 80.240 ;
        RECT 93.825 79.140 94.225 80.240 ;
        RECT 95.825 79.140 96.225 80.240 ;
        RECT 97.825 79.140 98.225 80.240 ;
        RECT 99.825 79.140 100.225 80.240 ;
        RECT 101.825 79.140 102.225 80.240 ;
        RECT 103.825 79.140 104.225 80.240 ;
        RECT 105.825 79.140 106.225 80.240 ;
        RECT 107.825 79.140 108.225 80.240 ;
        RECT 109.825 79.140 110.225 80.240 ;
        RECT 111.825 79.140 112.225 80.240 ;
        RECT 113.825 79.140 114.225 80.240 ;
        RECT 115.825 79.140 116.225 80.240 ;
        RECT 117.825 79.140 118.225 80.240 ;
        RECT 119.825 79.140 120.225 80.240 ;
        RECT 121.825 79.140 122.225 80.240 ;
        RECT 123.825 79.140 124.225 80.240 ;
        RECT 125.825 79.140 126.225 80.240 ;
        RECT 127.825 79.140 128.225 80.240 ;
        RECT 129.825 79.140 130.225 80.240 ;
        RECT 131.825 79.140 132.225 80.240 ;
        RECT 133.825 79.140 134.225 80.240 ;
        RECT 135.825 79.140 136.225 80.240 ;
        RECT 137.825 79.140 138.225 80.240 ;
        RECT 139.825 79.140 140.225 80.240 ;
        RECT 141.825 79.140 142.225 80.240 ;
        RECT 143.825 79.140 144.225 80.240 ;
        RECT 145.825 79.140 146.225 80.240 ;
        RECT 147.825 79.140 148.225 80.240 ;
        RECT 149.825 79.140 150.225 80.240 ;
        RECT 151.825 79.140 152.225 80.240 ;
        RECT 153.825 79.140 154.225 80.240 ;
        RECT 87.825 77.290 88.225 78.390 ;
        RECT 89.825 77.290 90.225 78.390 ;
        RECT 91.825 77.290 92.225 78.390 ;
        RECT 93.825 77.290 94.225 78.390 ;
        RECT 95.825 77.290 96.225 78.390 ;
        RECT 97.825 77.290 98.225 78.390 ;
        RECT 99.825 77.290 100.225 78.390 ;
        RECT 101.825 77.290 102.225 78.390 ;
        RECT 103.825 77.290 104.225 78.390 ;
        RECT 105.825 77.290 106.225 78.390 ;
        RECT 107.825 77.290 108.225 78.390 ;
        RECT 109.825 77.290 110.225 78.390 ;
        RECT 111.825 77.290 112.225 78.390 ;
        RECT 113.825 77.290 114.225 78.390 ;
        RECT 115.825 77.290 116.225 78.390 ;
        RECT 117.825 77.290 118.225 78.390 ;
        RECT 119.825 77.290 120.225 78.390 ;
        RECT 121.825 77.290 122.225 78.390 ;
        RECT 123.825 77.290 124.225 78.390 ;
        RECT 125.825 77.290 126.225 78.390 ;
        RECT 127.825 77.290 128.225 78.390 ;
        RECT 129.825 77.290 130.225 78.390 ;
        RECT 131.825 77.290 132.225 78.390 ;
        RECT 133.825 77.290 134.225 78.390 ;
        RECT 135.825 77.290 136.225 78.390 ;
        RECT 137.825 77.290 138.225 78.390 ;
        RECT 139.825 77.290 140.225 78.390 ;
        RECT 141.825 77.290 142.225 78.390 ;
        RECT 143.825 77.290 144.225 78.390 ;
        RECT 145.825 77.290 146.225 78.390 ;
        RECT 147.825 77.290 148.225 78.390 ;
        RECT 149.825 77.290 150.225 78.390 ;
        RECT 151.825 77.290 152.225 78.390 ;
        RECT 153.825 77.290 154.225 78.390 ;
        RECT 87.825 75.440 88.225 76.540 ;
        RECT 89.825 75.440 90.225 76.540 ;
        RECT 91.825 75.440 92.225 76.540 ;
        RECT 93.825 75.440 94.225 76.540 ;
        RECT 95.825 75.440 96.225 76.540 ;
        RECT 97.825 75.440 98.225 76.540 ;
        RECT 99.825 75.440 100.225 76.540 ;
        RECT 101.825 75.440 102.225 76.540 ;
        RECT 103.825 75.440 104.225 76.540 ;
        RECT 105.825 75.440 106.225 76.540 ;
        RECT 107.825 75.440 108.225 76.540 ;
        RECT 109.825 75.440 110.225 76.540 ;
        RECT 111.825 75.440 112.225 76.540 ;
        RECT 113.825 75.440 114.225 76.540 ;
        RECT 115.825 75.440 116.225 76.540 ;
        RECT 117.825 75.440 118.225 76.540 ;
        RECT 119.825 75.440 120.225 76.540 ;
        RECT 121.825 75.440 122.225 76.540 ;
        RECT 123.825 75.440 124.225 76.540 ;
        RECT 125.825 75.440 126.225 76.540 ;
        RECT 127.825 75.440 128.225 76.540 ;
        RECT 129.825 75.440 130.225 76.540 ;
        RECT 131.825 75.440 132.225 76.540 ;
        RECT 133.825 75.440 134.225 76.540 ;
        RECT 135.825 75.440 136.225 76.540 ;
        RECT 137.825 75.440 138.225 76.540 ;
        RECT 139.825 75.440 140.225 76.540 ;
        RECT 141.825 75.440 142.225 76.540 ;
        RECT 143.825 75.440 144.225 76.540 ;
        RECT 145.825 75.440 146.225 76.540 ;
        RECT 147.825 75.440 148.225 76.540 ;
        RECT 149.825 75.440 150.225 76.540 ;
        RECT 151.825 75.440 152.225 76.540 ;
        RECT 153.825 75.440 154.225 76.540 ;
        RECT 87.825 73.590 88.225 74.690 ;
        RECT 89.825 73.590 90.225 74.690 ;
        RECT 91.825 73.590 92.225 74.690 ;
        RECT 93.825 73.590 94.225 74.690 ;
        RECT 95.825 73.590 96.225 74.690 ;
        RECT 97.825 73.590 98.225 74.690 ;
        RECT 99.825 73.590 100.225 74.690 ;
        RECT 101.825 73.590 102.225 74.690 ;
        RECT 103.825 73.590 104.225 74.690 ;
        RECT 105.825 73.590 106.225 74.690 ;
        RECT 107.825 73.590 108.225 74.690 ;
        RECT 109.825 73.590 110.225 74.690 ;
        RECT 111.825 73.590 112.225 74.690 ;
        RECT 113.825 73.590 114.225 74.690 ;
        RECT 115.825 73.590 116.225 74.690 ;
        RECT 117.825 73.590 118.225 74.690 ;
        RECT 119.825 73.590 120.225 74.690 ;
        RECT 121.825 73.590 122.225 74.690 ;
        RECT 123.825 73.590 124.225 74.690 ;
        RECT 125.825 73.590 126.225 74.690 ;
        RECT 127.825 73.590 128.225 74.690 ;
        RECT 129.825 73.590 130.225 74.690 ;
        RECT 131.825 73.590 132.225 74.690 ;
        RECT 133.825 73.590 134.225 74.690 ;
        RECT 135.825 73.590 136.225 74.690 ;
        RECT 137.825 73.590 138.225 74.690 ;
        RECT 139.825 73.590 140.225 74.690 ;
        RECT 141.825 73.590 142.225 74.690 ;
        RECT 143.825 73.590 144.225 74.690 ;
        RECT 145.825 73.590 146.225 74.690 ;
        RECT 147.825 73.590 148.225 74.690 ;
        RECT 149.825 73.590 150.225 74.690 ;
        RECT 151.825 73.590 152.225 74.690 ;
        RECT 153.825 73.590 154.225 74.690 ;
        RECT 87.825 71.740 88.225 72.840 ;
        RECT 89.825 71.740 90.225 72.840 ;
        RECT 91.825 71.740 92.225 72.840 ;
        RECT 93.825 71.740 94.225 72.840 ;
        RECT 95.825 71.740 96.225 72.840 ;
        RECT 97.825 71.740 98.225 72.840 ;
        RECT 99.825 71.740 100.225 72.840 ;
        RECT 101.825 71.740 102.225 72.840 ;
        RECT 103.825 71.740 104.225 72.840 ;
        RECT 105.825 71.740 106.225 72.840 ;
        RECT 107.825 71.740 108.225 72.840 ;
        RECT 109.825 71.740 110.225 72.840 ;
        RECT 111.825 71.740 112.225 72.840 ;
        RECT 113.825 71.740 114.225 72.840 ;
        RECT 115.825 71.740 116.225 72.840 ;
        RECT 117.825 71.740 118.225 72.840 ;
        RECT 119.825 71.740 120.225 72.840 ;
        RECT 121.825 71.740 122.225 72.840 ;
        RECT 123.825 71.740 124.225 72.840 ;
        RECT 125.825 71.740 126.225 72.840 ;
        RECT 127.825 71.740 128.225 72.840 ;
        RECT 129.825 71.740 130.225 72.840 ;
        RECT 131.825 71.740 132.225 72.840 ;
        RECT 133.825 71.740 134.225 72.840 ;
        RECT 135.825 71.740 136.225 72.840 ;
        RECT 137.825 71.740 138.225 72.840 ;
        RECT 139.825 71.740 140.225 72.840 ;
        RECT 141.825 71.740 142.225 72.840 ;
        RECT 143.825 71.740 144.225 72.840 ;
        RECT 145.825 71.740 146.225 72.840 ;
        RECT 147.825 71.740 148.225 72.840 ;
        RECT 149.825 71.740 150.225 72.840 ;
        RECT 151.825 71.740 152.225 72.840 ;
        RECT 153.825 71.740 154.225 72.840 ;
        RECT 87.825 69.890 88.225 70.990 ;
        RECT 89.825 69.890 90.225 70.990 ;
        RECT 91.825 69.890 92.225 70.990 ;
        RECT 93.825 69.890 94.225 70.990 ;
        RECT 95.825 69.890 96.225 70.990 ;
        RECT 97.825 69.890 98.225 70.990 ;
        RECT 99.825 69.890 100.225 70.990 ;
        RECT 101.825 69.890 102.225 70.990 ;
        RECT 103.825 69.890 104.225 70.990 ;
        RECT 105.825 69.890 106.225 70.990 ;
        RECT 107.825 69.890 108.225 70.990 ;
        RECT 109.825 69.890 110.225 70.990 ;
        RECT 111.825 69.890 112.225 70.990 ;
        RECT 113.825 69.890 114.225 70.990 ;
        RECT 115.825 69.890 116.225 70.990 ;
        RECT 117.825 69.890 118.225 70.990 ;
        RECT 119.825 69.890 120.225 70.990 ;
        RECT 121.825 69.890 122.225 70.990 ;
        RECT 123.825 69.890 124.225 70.990 ;
        RECT 125.825 69.890 126.225 70.990 ;
        RECT 127.825 69.890 128.225 70.990 ;
        RECT 129.825 69.890 130.225 70.990 ;
        RECT 131.825 69.890 132.225 70.990 ;
        RECT 133.825 69.890 134.225 70.990 ;
        RECT 135.825 69.890 136.225 70.990 ;
        RECT 137.825 69.890 138.225 70.990 ;
        RECT 139.825 69.890 140.225 70.990 ;
        RECT 141.825 69.890 142.225 70.990 ;
        RECT 143.825 69.890 144.225 70.990 ;
        RECT 145.825 69.890 146.225 70.990 ;
        RECT 147.825 69.890 148.225 70.990 ;
        RECT 149.825 69.890 150.225 70.990 ;
        RECT 151.825 69.890 152.225 70.990 ;
        RECT 153.825 69.890 154.225 70.990 ;
        RECT 87.825 68.040 88.225 69.140 ;
        RECT 89.825 68.040 90.225 69.140 ;
        RECT 91.825 68.040 92.225 69.140 ;
        RECT 93.825 68.040 94.225 69.140 ;
        RECT 95.825 68.040 96.225 69.140 ;
        RECT 97.825 68.040 98.225 69.140 ;
        RECT 99.825 68.040 100.225 69.140 ;
        RECT 101.825 68.040 102.225 69.140 ;
        RECT 103.825 68.040 104.225 69.140 ;
        RECT 105.825 68.040 106.225 69.140 ;
        RECT 107.825 68.040 108.225 69.140 ;
        RECT 109.825 68.040 110.225 69.140 ;
        RECT 111.825 68.040 112.225 69.140 ;
        RECT 113.825 68.040 114.225 69.140 ;
        RECT 115.825 68.040 116.225 69.140 ;
        RECT 117.825 68.040 118.225 69.140 ;
        RECT 119.825 68.040 120.225 69.140 ;
        RECT 121.825 68.040 122.225 69.140 ;
        RECT 123.825 68.040 124.225 69.140 ;
        RECT 125.825 68.040 126.225 69.140 ;
        RECT 127.825 68.040 128.225 69.140 ;
        RECT 129.825 68.040 130.225 69.140 ;
        RECT 131.825 68.040 132.225 69.140 ;
        RECT 133.825 68.040 134.225 69.140 ;
        RECT 135.825 68.040 136.225 69.140 ;
        RECT 137.825 68.040 138.225 69.140 ;
        RECT 139.825 68.040 140.225 69.140 ;
        RECT 141.825 68.040 142.225 69.140 ;
        RECT 143.825 68.040 144.225 69.140 ;
        RECT 145.825 68.040 146.225 69.140 ;
        RECT 147.825 68.040 148.225 69.140 ;
        RECT 149.825 68.040 150.225 69.140 ;
        RECT 151.825 68.040 152.225 69.140 ;
        RECT 153.825 68.040 154.225 69.140 ;
        RECT 87.825 66.190 88.225 67.290 ;
        RECT 89.825 66.190 90.225 67.290 ;
        RECT 91.825 66.190 92.225 67.290 ;
        RECT 93.825 66.190 94.225 67.290 ;
        RECT 95.825 66.190 96.225 67.290 ;
        RECT 97.825 66.190 98.225 67.290 ;
        RECT 99.825 66.190 100.225 67.290 ;
        RECT 101.825 66.190 102.225 67.290 ;
        RECT 103.825 66.190 104.225 67.290 ;
        RECT 105.825 66.190 106.225 67.290 ;
        RECT 107.825 66.190 108.225 67.290 ;
        RECT 109.825 66.190 110.225 67.290 ;
        RECT 111.825 66.190 112.225 67.290 ;
        RECT 113.825 66.190 114.225 67.290 ;
        RECT 115.825 66.190 116.225 67.290 ;
        RECT 117.825 66.190 118.225 67.290 ;
        RECT 119.825 66.190 120.225 67.290 ;
        RECT 121.825 66.190 122.225 67.290 ;
        RECT 123.825 66.190 124.225 67.290 ;
        RECT 125.825 66.190 126.225 67.290 ;
        RECT 127.825 66.190 128.225 67.290 ;
        RECT 129.825 66.190 130.225 67.290 ;
        RECT 131.825 66.190 132.225 67.290 ;
        RECT 133.825 66.190 134.225 67.290 ;
        RECT 135.825 66.190 136.225 67.290 ;
        RECT 137.825 66.190 138.225 67.290 ;
        RECT 139.825 66.190 140.225 67.290 ;
        RECT 141.825 66.190 142.225 67.290 ;
        RECT 143.825 66.190 144.225 67.290 ;
        RECT 145.825 66.190 146.225 67.290 ;
        RECT 147.825 66.190 148.225 67.290 ;
        RECT 149.825 66.190 150.225 67.290 ;
        RECT 151.825 66.190 152.225 67.290 ;
        RECT 153.825 66.190 154.225 67.290 ;
        RECT 87.825 64.340 88.225 65.440 ;
        RECT 89.825 64.340 90.225 65.440 ;
        RECT 91.825 64.340 92.225 65.440 ;
        RECT 93.825 64.340 94.225 65.440 ;
        RECT 95.825 64.340 96.225 65.440 ;
        RECT 97.825 64.340 98.225 65.440 ;
        RECT 99.825 64.340 100.225 65.440 ;
        RECT 101.825 64.340 102.225 65.440 ;
        RECT 103.825 64.340 104.225 65.440 ;
        RECT 105.825 64.340 106.225 65.440 ;
        RECT 107.825 64.340 108.225 65.440 ;
        RECT 109.825 64.340 110.225 65.440 ;
        RECT 111.825 64.340 112.225 65.440 ;
        RECT 113.825 64.340 114.225 65.440 ;
        RECT 115.825 64.340 116.225 65.440 ;
        RECT 117.825 64.340 118.225 65.440 ;
        RECT 119.825 64.340 120.225 65.440 ;
        RECT 121.825 64.340 122.225 65.440 ;
        RECT 123.825 64.340 124.225 65.440 ;
        RECT 125.825 64.340 126.225 65.440 ;
        RECT 127.825 64.340 128.225 65.440 ;
        RECT 129.825 64.340 130.225 65.440 ;
        RECT 131.825 64.340 132.225 65.440 ;
        RECT 133.825 64.340 134.225 65.440 ;
        RECT 135.825 64.340 136.225 65.440 ;
        RECT 137.825 64.340 138.225 65.440 ;
        RECT 139.825 64.340 140.225 65.440 ;
        RECT 141.825 64.340 142.225 65.440 ;
        RECT 143.825 64.340 144.225 65.440 ;
        RECT 145.825 64.340 146.225 65.440 ;
        RECT 147.825 64.340 148.225 65.440 ;
        RECT 149.825 64.340 150.225 65.440 ;
        RECT 151.825 64.340 152.225 65.440 ;
        RECT 153.825 64.340 154.225 65.440 ;
        RECT 87.825 62.490 88.225 63.590 ;
        RECT 89.825 62.490 90.225 63.590 ;
        RECT 91.825 62.490 92.225 63.590 ;
        RECT 93.825 62.490 94.225 63.590 ;
        RECT 95.825 62.490 96.225 63.590 ;
        RECT 97.825 62.490 98.225 63.590 ;
        RECT 99.825 62.490 100.225 63.590 ;
        RECT 101.825 62.490 102.225 63.590 ;
        RECT 103.825 62.490 104.225 63.590 ;
        RECT 105.825 62.490 106.225 63.590 ;
        RECT 107.825 62.490 108.225 63.590 ;
        RECT 109.825 62.490 110.225 63.590 ;
        RECT 111.825 62.490 112.225 63.590 ;
        RECT 113.825 62.490 114.225 63.590 ;
        RECT 115.825 62.490 116.225 63.590 ;
        RECT 117.825 62.490 118.225 63.590 ;
        RECT 119.825 62.490 120.225 63.590 ;
        RECT 121.825 62.490 122.225 63.590 ;
        RECT 123.825 62.490 124.225 63.590 ;
        RECT 125.825 62.490 126.225 63.590 ;
        RECT 127.825 62.490 128.225 63.590 ;
        RECT 129.825 62.490 130.225 63.590 ;
        RECT 131.825 62.490 132.225 63.590 ;
        RECT 133.825 62.490 134.225 63.590 ;
        RECT 135.825 62.490 136.225 63.590 ;
        RECT 137.825 62.490 138.225 63.590 ;
        RECT 139.825 62.490 140.225 63.590 ;
        RECT 141.825 62.490 142.225 63.590 ;
        RECT 143.825 62.490 144.225 63.590 ;
        RECT 145.825 62.490 146.225 63.590 ;
        RECT 147.825 62.490 148.225 63.590 ;
        RECT 149.825 62.490 150.225 63.590 ;
        RECT 151.825 62.490 152.225 63.590 ;
        RECT 153.825 62.490 154.225 63.590 ;
        RECT 87.825 60.640 88.225 61.740 ;
        RECT 89.825 60.640 90.225 61.740 ;
        RECT 91.825 60.640 92.225 61.740 ;
        RECT 93.825 60.640 94.225 61.740 ;
        RECT 95.825 60.640 96.225 61.740 ;
        RECT 97.825 60.640 98.225 61.740 ;
        RECT 99.825 60.640 100.225 61.740 ;
        RECT 101.825 60.640 102.225 61.740 ;
        RECT 103.825 60.640 104.225 61.740 ;
        RECT 105.825 60.640 106.225 61.740 ;
        RECT 107.825 60.640 108.225 61.740 ;
        RECT 109.825 60.640 110.225 61.740 ;
        RECT 111.825 60.640 112.225 61.740 ;
        RECT 113.825 60.640 114.225 61.740 ;
        RECT 115.825 60.640 116.225 61.740 ;
        RECT 117.825 60.640 118.225 61.740 ;
        RECT 119.825 60.640 120.225 61.740 ;
        RECT 121.825 60.640 122.225 61.740 ;
        RECT 123.825 60.640 124.225 61.740 ;
        RECT 125.825 60.640 126.225 61.740 ;
        RECT 127.825 60.640 128.225 61.740 ;
        RECT 129.825 60.640 130.225 61.740 ;
        RECT 131.825 60.640 132.225 61.740 ;
        RECT 133.825 60.640 134.225 61.740 ;
        RECT 135.825 60.640 136.225 61.740 ;
        RECT 137.825 60.640 138.225 61.740 ;
        RECT 139.825 60.640 140.225 61.740 ;
        RECT 141.825 60.640 142.225 61.740 ;
        RECT 143.825 60.640 144.225 61.740 ;
        RECT 145.825 60.640 146.225 61.740 ;
        RECT 147.825 60.640 148.225 61.740 ;
        RECT 149.825 60.640 150.225 61.740 ;
        RECT 151.825 60.640 152.225 61.740 ;
        RECT 153.825 60.640 154.225 61.740 ;
        RECT 87.825 58.790 88.225 59.890 ;
        RECT 89.825 58.790 90.225 59.890 ;
        RECT 91.825 58.790 92.225 59.890 ;
        RECT 93.825 58.790 94.225 59.890 ;
        RECT 95.825 58.790 96.225 59.890 ;
        RECT 97.825 58.790 98.225 59.890 ;
        RECT 99.825 58.790 100.225 59.890 ;
        RECT 101.825 58.790 102.225 59.890 ;
        RECT 103.825 58.790 104.225 59.890 ;
        RECT 105.825 58.790 106.225 59.890 ;
        RECT 107.825 58.790 108.225 59.890 ;
        RECT 109.825 58.790 110.225 59.890 ;
        RECT 111.825 58.790 112.225 59.890 ;
        RECT 113.825 58.790 114.225 59.890 ;
        RECT 115.825 58.790 116.225 59.890 ;
        RECT 117.825 58.790 118.225 59.890 ;
        RECT 119.825 58.790 120.225 59.890 ;
        RECT 121.825 58.790 122.225 59.890 ;
        RECT 123.825 58.790 124.225 59.890 ;
        RECT 125.825 58.790 126.225 59.890 ;
        RECT 127.825 58.790 128.225 59.890 ;
        RECT 129.825 58.790 130.225 59.890 ;
        RECT 131.825 58.790 132.225 59.890 ;
        RECT 133.825 58.790 134.225 59.890 ;
        RECT 135.825 58.790 136.225 59.890 ;
        RECT 137.825 58.790 138.225 59.890 ;
        RECT 139.825 58.790 140.225 59.890 ;
        RECT 141.825 58.790 142.225 59.890 ;
        RECT 143.825 58.790 144.225 59.890 ;
        RECT 145.825 58.790 146.225 59.890 ;
        RECT 147.825 58.790 148.225 59.890 ;
        RECT 149.825 58.790 150.225 59.890 ;
        RECT 151.825 58.790 152.225 59.890 ;
        RECT 153.825 58.790 154.225 59.890 ;
        RECT 87.825 56.940 88.225 58.040 ;
        RECT 89.825 56.940 90.225 58.040 ;
        RECT 91.825 56.940 92.225 58.040 ;
        RECT 93.825 56.940 94.225 58.040 ;
        RECT 95.825 56.940 96.225 58.040 ;
        RECT 97.825 56.940 98.225 58.040 ;
        RECT 99.825 56.940 100.225 58.040 ;
        RECT 101.825 56.940 102.225 58.040 ;
        RECT 103.825 56.940 104.225 58.040 ;
        RECT 105.825 56.940 106.225 58.040 ;
        RECT 107.825 56.940 108.225 58.040 ;
        RECT 109.825 56.940 110.225 58.040 ;
        RECT 111.825 56.940 112.225 58.040 ;
        RECT 113.825 56.940 114.225 58.040 ;
        RECT 115.825 56.940 116.225 58.040 ;
        RECT 117.825 56.940 118.225 58.040 ;
        RECT 119.825 56.940 120.225 58.040 ;
        RECT 121.825 56.940 122.225 58.040 ;
        RECT 123.825 56.940 124.225 58.040 ;
        RECT 125.825 56.940 126.225 58.040 ;
        RECT 127.825 56.940 128.225 58.040 ;
        RECT 129.825 56.940 130.225 58.040 ;
        RECT 131.825 56.940 132.225 58.040 ;
        RECT 133.825 56.940 134.225 58.040 ;
        RECT 135.825 56.940 136.225 58.040 ;
        RECT 137.825 56.940 138.225 58.040 ;
        RECT 139.825 56.940 140.225 58.040 ;
        RECT 141.825 56.940 142.225 58.040 ;
        RECT 143.825 56.940 144.225 58.040 ;
        RECT 145.825 56.940 146.225 58.040 ;
        RECT 147.825 56.940 148.225 58.040 ;
        RECT 149.825 56.940 150.225 58.040 ;
        RECT 151.825 56.940 152.225 58.040 ;
        RECT 153.825 56.940 154.225 58.040 ;
        RECT 87.825 55.090 88.225 56.190 ;
        RECT 89.825 55.090 90.225 56.190 ;
        RECT 91.825 55.090 92.225 56.190 ;
        RECT 93.825 55.090 94.225 56.190 ;
        RECT 95.825 55.090 96.225 56.190 ;
        RECT 97.825 55.090 98.225 56.190 ;
        RECT 99.825 55.090 100.225 56.190 ;
        RECT 101.825 55.090 102.225 56.190 ;
        RECT 103.825 55.090 104.225 56.190 ;
        RECT 105.825 55.090 106.225 56.190 ;
        RECT 107.825 55.090 108.225 56.190 ;
        RECT 109.825 55.090 110.225 56.190 ;
        RECT 111.825 55.090 112.225 56.190 ;
        RECT 113.825 55.090 114.225 56.190 ;
        RECT 115.825 55.090 116.225 56.190 ;
        RECT 117.825 55.090 118.225 56.190 ;
        RECT 119.825 55.090 120.225 56.190 ;
        RECT 121.825 55.090 122.225 56.190 ;
        RECT 123.825 55.090 124.225 56.190 ;
        RECT 125.825 55.090 126.225 56.190 ;
        RECT 127.825 55.090 128.225 56.190 ;
        RECT 129.825 55.090 130.225 56.190 ;
        RECT 131.825 55.090 132.225 56.190 ;
        RECT 133.825 55.090 134.225 56.190 ;
        RECT 135.825 55.090 136.225 56.190 ;
        RECT 137.825 55.090 138.225 56.190 ;
        RECT 139.825 55.090 140.225 56.190 ;
        RECT 141.825 55.090 142.225 56.190 ;
        RECT 143.825 55.090 144.225 56.190 ;
        RECT 145.825 55.090 146.225 56.190 ;
        RECT 147.825 55.090 148.225 56.190 ;
        RECT 149.825 55.090 150.225 56.190 ;
        RECT 151.825 55.090 152.225 56.190 ;
        RECT 153.825 55.090 154.225 56.190 ;
        RECT 87.825 53.240 88.225 54.340 ;
        RECT 89.825 53.240 90.225 54.340 ;
        RECT 91.825 53.240 92.225 54.340 ;
        RECT 93.825 53.240 94.225 54.340 ;
        RECT 95.825 53.240 96.225 54.340 ;
        RECT 97.825 53.240 98.225 54.340 ;
        RECT 99.825 53.240 100.225 54.340 ;
        RECT 101.825 53.240 102.225 54.340 ;
        RECT 103.825 53.240 104.225 54.340 ;
        RECT 105.825 53.240 106.225 54.340 ;
        RECT 107.825 53.240 108.225 54.340 ;
        RECT 109.825 53.240 110.225 54.340 ;
        RECT 111.825 53.240 112.225 54.340 ;
        RECT 113.825 53.240 114.225 54.340 ;
        RECT 115.825 53.240 116.225 54.340 ;
        RECT 117.825 53.240 118.225 54.340 ;
        RECT 119.825 53.240 120.225 54.340 ;
        RECT 121.825 53.240 122.225 54.340 ;
        RECT 123.825 53.240 124.225 54.340 ;
        RECT 125.825 53.240 126.225 54.340 ;
        RECT 127.825 53.240 128.225 54.340 ;
        RECT 129.825 53.240 130.225 54.340 ;
        RECT 131.825 53.240 132.225 54.340 ;
        RECT 133.825 53.240 134.225 54.340 ;
        RECT 135.825 53.240 136.225 54.340 ;
        RECT 137.825 53.240 138.225 54.340 ;
        RECT 139.825 53.240 140.225 54.340 ;
        RECT 141.825 53.240 142.225 54.340 ;
        RECT 143.825 53.240 144.225 54.340 ;
        RECT 145.825 53.240 146.225 54.340 ;
        RECT 147.825 53.240 148.225 54.340 ;
        RECT 149.825 53.240 150.225 54.340 ;
        RECT 151.825 53.240 152.225 54.340 ;
        RECT 153.825 53.240 154.225 54.340 ;
        RECT 87.825 51.390 88.225 52.490 ;
        RECT 89.825 51.390 90.225 52.490 ;
        RECT 91.825 51.390 92.225 52.490 ;
        RECT 93.825 51.390 94.225 52.490 ;
        RECT 95.825 51.390 96.225 52.490 ;
        RECT 97.825 51.390 98.225 52.490 ;
        RECT 99.825 51.390 100.225 52.490 ;
        RECT 101.825 51.390 102.225 52.490 ;
        RECT 103.825 51.390 104.225 52.490 ;
        RECT 105.825 51.390 106.225 52.490 ;
        RECT 107.825 51.390 108.225 52.490 ;
        RECT 109.825 51.390 110.225 52.490 ;
        RECT 111.825 51.390 112.225 52.490 ;
        RECT 113.825 51.390 114.225 52.490 ;
        RECT 115.825 51.390 116.225 52.490 ;
        RECT 117.825 51.390 118.225 52.490 ;
        RECT 119.825 51.390 120.225 52.490 ;
        RECT 121.825 51.390 122.225 52.490 ;
        RECT 123.825 51.390 124.225 52.490 ;
        RECT 125.825 51.390 126.225 52.490 ;
        RECT 127.825 51.390 128.225 52.490 ;
        RECT 129.825 51.390 130.225 52.490 ;
        RECT 131.825 51.390 132.225 52.490 ;
        RECT 133.825 51.390 134.225 52.490 ;
        RECT 135.825 51.390 136.225 52.490 ;
        RECT 137.825 51.390 138.225 52.490 ;
        RECT 139.825 51.390 140.225 52.490 ;
        RECT 141.825 51.390 142.225 52.490 ;
        RECT 143.825 51.390 144.225 52.490 ;
        RECT 145.825 51.390 146.225 52.490 ;
        RECT 147.825 51.390 148.225 52.490 ;
        RECT 149.825 51.390 150.225 52.490 ;
        RECT 151.825 51.390 152.225 52.490 ;
        RECT 153.825 51.390 154.225 52.490 ;
        RECT 87.825 49.540 88.225 50.640 ;
        RECT 89.825 49.540 90.225 50.640 ;
        RECT 91.825 49.540 92.225 50.640 ;
        RECT 93.825 49.540 94.225 50.640 ;
        RECT 95.825 49.540 96.225 50.640 ;
        RECT 97.825 49.540 98.225 50.640 ;
        RECT 99.825 49.540 100.225 50.640 ;
        RECT 101.825 49.540 102.225 50.640 ;
        RECT 103.825 49.540 104.225 50.640 ;
        RECT 105.825 49.540 106.225 50.640 ;
        RECT 107.825 49.540 108.225 50.640 ;
        RECT 109.825 49.540 110.225 50.640 ;
        RECT 111.825 49.540 112.225 50.640 ;
        RECT 113.825 49.540 114.225 50.640 ;
        RECT 115.825 49.540 116.225 50.640 ;
        RECT 117.825 49.540 118.225 50.640 ;
        RECT 119.825 49.540 120.225 50.640 ;
        RECT 121.825 49.540 122.225 50.640 ;
        RECT 123.825 49.540 124.225 50.640 ;
        RECT 125.825 49.540 126.225 50.640 ;
        RECT 127.825 49.540 128.225 50.640 ;
        RECT 129.825 49.540 130.225 50.640 ;
        RECT 131.825 49.540 132.225 50.640 ;
        RECT 133.825 49.540 134.225 50.640 ;
        RECT 135.825 49.540 136.225 50.640 ;
        RECT 137.825 49.540 138.225 50.640 ;
        RECT 139.825 49.540 140.225 50.640 ;
        RECT 141.825 49.540 142.225 50.640 ;
        RECT 143.825 49.540 144.225 50.640 ;
        RECT 145.825 49.540 146.225 50.640 ;
        RECT 147.825 49.540 148.225 50.640 ;
        RECT 149.825 49.540 150.225 50.640 ;
        RECT 151.825 49.540 152.225 50.640 ;
        RECT 153.825 49.540 154.225 50.640 ;
        RECT 87.825 47.690 88.225 48.790 ;
        RECT 89.825 47.690 90.225 48.790 ;
        RECT 91.825 47.690 92.225 48.790 ;
        RECT 93.825 47.690 94.225 48.790 ;
        RECT 95.825 47.690 96.225 48.790 ;
        RECT 97.825 47.690 98.225 48.790 ;
        RECT 99.825 47.690 100.225 48.790 ;
        RECT 101.825 47.690 102.225 48.790 ;
        RECT 103.825 47.690 104.225 48.790 ;
        RECT 105.825 47.690 106.225 48.790 ;
        RECT 107.825 47.690 108.225 48.790 ;
        RECT 109.825 47.690 110.225 48.790 ;
        RECT 111.825 47.690 112.225 48.790 ;
        RECT 113.825 47.690 114.225 48.790 ;
        RECT 115.825 47.690 116.225 48.790 ;
        RECT 117.825 47.690 118.225 48.790 ;
        RECT 119.825 47.690 120.225 48.790 ;
        RECT 121.825 47.690 122.225 48.790 ;
        RECT 123.825 47.690 124.225 48.790 ;
        RECT 125.825 47.690 126.225 48.790 ;
        RECT 127.825 47.690 128.225 48.790 ;
        RECT 129.825 47.690 130.225 48.790 ;
        RECT 131.825 47.690 132.225 48.790 ;
        RECT 133.825 47.690 134.225 48.790 ;
        RECT 135.825 47.690 136.225 48.790 ;
        RECT 137.825 47.690 138.225 48.790 ;
        RECT 139.825 47.690 140.225 48.790 ;
        RECT 141.825 47.690 142.225 48.790 ;
        RECT 143.825 47.690 144.225 48.790 ;
        RECT 145.825 47.690 146.225 48.790 ;
        RECT 147.825 47.690 148.225 48.790 ;
        RECT 149.825 47.690 150.225 48.790 ;
        RECT 151.825 47.690 152.225 48.790 ;
        RECT 153.825 47.690 154.225 48.790 ;
        RECT 87.825 45.840 88.225 46.940 ;
        RECT 89.825 45.840 90.225 46.940 ;
        RECT 91.825 45.840 92.225 46.940 ;
        RECT 93.825 45.840 94.225 46.940 ;
        RECT 95.825 45.840 96.225 46.940 ;
        RECT 97.825 45.840 98.225 46.940 ;
        RECT 99.825 45.840 100.225 46.940 ;
        RECT 101.825 45.840 102.225 46.940 ;
        RECT 103.825 45.840 104.225 46.940 ;
        RECT 105.825 45.840 106.225 46.940 ;
        RECT 107.825 45.840 108.225 46.940 ;
        RECT 109.825 45.840 110.225 46.940 ;
        RECT 111.825 45.840 112.225 46.940 ;
        RECT 113.825 45.840 114.225 46.940 ;
        RECT 115.825 45.840 116.225 46.940 ;
        RECT 117.825 45.840 118.225 46.940 ;
        RECT 119.825 45.840 120.225 46.940 ;
        RECT 121.825 45.840 122.225 46.940 ;
        RECT 123.825 45.840 124.225 46.940 ;
        RECT 125.825 45.840 126.225 46.940 ;
        RECT 127.825 45.840 128.225 46.940 ;
        RECT 129.825 45.840 130.225 46.940 ;
        RECT 131.825 45.840 132.225 46.940 ;
        RECT 133.825 45.840 134.225 46.940 ;
        RECT 135.825 45.840 136.225 46.940 ;
        RECT 137.825 45.840 138.225 46.940 ;
        RECT 139.825 45.840 140.225 46.940 ;
        RECT 141.825 45.840 142.225 46.940 ;
        RECT 143.825 45.840 144.225 46.940 ;
        RECT 145.825 45.840 146.225 46.940 ;
        RECT 147.825 45.840 148.225 46.940 ;
        RECT 149.825 45.840 150.225 46.940 ;
        RECT 151.825 45.840 152.225 46.940 ;
        RECT 153.825 45.840 154.225 46.940 ;
        RECT 87.825 43.990 88.225 45.090 ;
        RECT 89.825 43.990 90.225 45.090 ;
        RECT 91.825 43.990 92.225 45.090 ;
        RECT 93.825 43.990 94.225 45.090 ;
        RECT 95.825 43.990 96.225 45.090 ;
        RECT 97.825 43.990 98.225 45.090 ;
        RECT 99.825 43.990 100.225 45.090 ;
        RECT 101.825 43.990 102.225 45.090 ;
        RECT 103.825 43.990 104.225 45.090 ;
        RECT 105.825 43.990 106.225 45.090 ;
        RECT 107.825 43.990 108.225 45.090 ;
        RECT 109.825 43.990 110.225 45.090 ;
        RECT 111.825 43.990 112.225 45.090 ;
        RECT 113.825 43.990 114.225 45.090 ;
        RECT 115.825 43.990 116.225 45.090 ;
        RECT 117.825 43.990 118.225 45.090 ;
        RECT 119.825 43.990 120.225 45.090 ;
        RECT 121.825 43.990 122.225 45.090 ;
        RECT 123.825 43.990 124.225 45.090 ;
        RECT 125.825 43.990 126.225 45.090 ;
        RECT 127.825 43.990 128.225 45.090 ;
        RECT 129.825 43.990 130.225 45.090 ;
        RECT 131.825 43.990 132.225 45.090 ;
        RECT 133.825 43.990 134.225 45.090 ;
        RECT 135.825 43.990 136.225 45.090 ;
        RECT 137.825 43.990 138.225 45.090 ;
        RECT 139.825 43.990 140.225 45.090 ;
        RECT 141.825 43.990 142.225 45.090 ;
        RECT 143.825 43.990 144.225 45.090 ;
        RECT 145.825 43.990 146.225 45.090 ;
        RECT 147.825 43.990 148.225 45.090 ;
        RECT 149.825 43.990 150.225 45.090 ;
        RECT 151.825 43.990 152.225 45.090 ;
        RECT 153.825 43.990 154.225 45.090 ;
        RECT 87.825 42.140 88.225 43.240 ;
        RECT 89.825 42.140 90.225 43.240 ;
        RECT 91.825 42.140 92.225 43.240 ;
        RECT 93.825 42.140 94.225 43.240 ;
        RECT 95.825 42.140 96.225 43.240 ;
        RECT 97.825 42.140 98.225 43.240 ;
        RECT 99.825 42.140 100.225 43.240 ;
        RECT 101.825 42.140 102.225 43.240 ;
        RECT 103.825 42.140 104.225 43.240 ;
        RECT 105.825 42.140 106.225 43.240 ;
        RECT 107.825 42.140 108.225 43.240 ;
        RECT 109.825 42.140 110.225 43.240 ;
        RECT 111.825 42.140 112.225 43.240 ;
        RECT 113.825 42.140 114.225 43.240 ;
        RECT 115.825 42.140 116.225 43.240 ;
        RECT 117.825 42.140 118.225 43.240 ;
        RECT 119.825 42.140 120.225 43.240 ;
        RECT 121.825 42.140 122.225 43.240 ;
        RECT 123.825 42.140 124.225 43.240 ;
        RECT 125.825 42.140 126.225 43.240 ;
        RECT 127.825 42.140 128.225 43.240 ;
        RECT 129.825 42.140 130.225 43.240 ;
        RECT 131.825 42.140 132.225 43.240 ;
        RECT 133.825 42.140 134.225 43.240 ;
        RECT 135.825 42.140 136.225 43.240 ;
        RECT 137.825 42.140 138.225 43.240 ;
        RECT 139.825 42.140 140.225 43.240 ;
        RECT 141.825 42.140 142.225 43.240 ;
        RECT 143.825 42.140 144.225 43.240 ;
        RECT 145.825 42.140 146.225 43.240 ;
        RECT 147.825 42.140 148.225 43.240 ;
        RECT 149.825 42.140 150.225 43.240 ;
        RECT 151.825 42.140 152.225 43.240 ;
        RECT 153.825 42.140 154.225 43.240 ;
        RECT 87.825 40.290 88.225 41.390 ;
        RECT 89.825 40.290 90.225 41.390 ;
        RECT 91.825 40.290 92.225 41.390 ;
        RECT 93.825 40.290 94.225 41.390 ;
        RECT 95.825 40.290 96.225 41.390 ;
        RECT 97.825 40.290 98.225 41.390 ;
        RECT 99.825 40.290 100.225 41.390 ;
        RECT 101.825 40.290 102.225 41.390 ;
        RECT 103.825 40.290 104.225 41.390 ;
        RECT 105.825 40.290 106.225 41.390 ;
        RECT 107.825 40.290 108.225 41.390 ;
        RECT 109.825 40.290 110.225 41.390 ;
        RECT 111.825 40.290 112.225 41.390 ;
        RECT 113.825 40.290 114.225 41.390 ;
        RECT 115.825 40.290 116.225 41.390 ;
        RECT 117.825 40.290 118.225 41.390 ;
        RECT 119.825 40.290 120.225 41.390 ;
        RECT 121.825 40.290 122.225 41.390 ;
        RECT 123.825 40.290 124.225 41.390 ;
        RECT 125.825 40.290 126.225 41.390 ;
        RECT 127.825 40.290 128.225 41.390 ;
        RECT 129.825 40.290 130.225 41.390 ;
        RECT 131.825 40.290 132.225 41.390 ;
        RECT 133.825 40.290 134.225 41.390 ;
        RECT 135.825 40.290 136.225 41.390 ;
        RECT 137.825 40.290 138.225 41.390 ;
        RECT 139.825 40.290 140.225 41.390 ;
        RECT 141.825 40.290 142.225 41.390 ;
        RECT 143.825 40.290 144.225 41.390 ;
        RECT 145.825 40.290 146.225 41.390 ;
        RECT 147.825 40.290 148.225 41.390 ;
        RECT 149.825 40.290 150.225 41.390 ;
        RECT 151.825 40.290 152.225 41.390 ;
        RECT 153.825 40.290 154.225 41.390 ;
        RECT 87.825 38.440 88.225 39.540 ;
        RECT 89.825 38.440 90.225 39.540 ;
        RECT 91.825 38.440 92.225 39.540 ;
        RECT 93.825 38.440 94.225 39.540 ;
        RECT 95.825 38.440 96.225 39.540 ;
        RECT 97.825 38.440 98.225 39.540 ;
        RECT 99.825 38.440 100.225 39.540 ;
        RECT 101.825 38.440 102.225 39.540 ;
        RECT 103.825 38.440 104.225 39.540 ;
        RECT 105.825 38.440 106.225 39.540 ;
        RECT 107.825 38.440 108.225 39.540 ;
        RECT 109.825 38.440 110.225 39.540 ;
        RECT 111.825 38.440 112.225 39.540 ;
        RECT 113.825 38.440 114.225 39.540 ;
        RECT 115.825 38.440 116.225 39.540 ;
        RECT 117.825 38.440 118.225 39.540 ;
        RECT 119.825 38.440 120.225 39.540 ;
        RECT 121.825 38.440 122.225 39.540 ;
        RECT 123.825 38.440 124.225 39.540 ;
        RECT 125.825 38.440 126.225 39.540 ;
        RECT 127.825 38.440 128.225 39.540 ;
        RECT 129.825 38.440 130.225 39.540 ;
        RECT 131.825 38.440 132.225 39.540 ;
        RECT 133.825 38.440 134.225 39.540 ;
        RECT 135.825 38.440 136.225 39.540 ;
        RECT 137.825 38.440 138.225 39.540 ;
        RECT 139.825 38.440 140.225 39.540 ;
        RECT 141.825 38.440 142.225 39.540 ;
        RECT 143.825 38.440 144.225 39.540 ;
        RECT 145.825 38.440 146.225 39.540 ;
        RECT 147.825 38.440 148.225 39.540 ;
        RECT 149.825 38.440 150.225 39.540 ;
        RECT 151.825 38.440 152.225 39.540 ;
        RECT 153.825 38.440 154.225 39.540 ;
        RECT 87.825 36.590 88.225 37.690 ;
        RECT 89.825 36.590 90.225 37.690 ;
        RECT 91.825 36.590 92.225 37.690 ;
        RECT 93.825 36.590 94.225 37.690 ;
        RECT 95.825 36.590 96.225 37.690 ;
        RECT 97.825 36.590 98.225 37.690 ;
        RECT 99.825 36.590 100.225 37.690 ;
        RECT 101.825 36.590 102.225 37.690 ;
        RECT 103.825 36.590 104.225 37.690 ;
        RECT 105.825 36.590 106.225 37.690 ;
        RECT 107.825 36.590 108.225 37.690 ;
        RECT 109.825 36.590 110.225 37.690 ;
        RECT 111.825 36.590 112.225 37.690 ;
        RECT 113.825 36.590 114.225 37.690 ;
        RECT 115.825 36.590 116.225 37.690 ;
        RECT 117.825 36.590 118.225 37.690 ;
        RECT 119.825 36.590 120.225 37.690 ;
        RECT 121.825 36.590 122.225 37.690 ;
        RECT 123.825 36.590 124.225 37.690 ;
        RECT 125.825 36.590 126.225 37.690 ;
        RECT 127.825 36.590 128.225 37.690 ;
        RECT 129.825 36.590 130.225 37.690 ;
        RECT 131.825 36.590 132.225 37.690 ;
        RECT 133.825 36.590 134.225 37.690 ;
        RECT 135.825 36.590 136.225 37.690 ;
        RECT 137.825 36.590 138.225 37.690 ;
        RECT 139.825 36.590 140.225 37.690 ;
        RECT 141.825 36.590 142.225 37.690 ;
        RECT 143.825 36.590 144.225 37.690 ;
        RECT 145.825 36.590 146.225 37.690 ;
        RECT 147.825 36.590 148.225 37.690 ;
        RECT 149.825 36.590 150.225 37.690 ;
        RECT 151.825 36.590 152.225 37.690 ;
        RECT 153.825 36.590 154.225 37.690 ;
        RECT 87.825 34.740 88.225 35.840 ;
        RECT 89.825 34.740 90.225 35.840 ;
        RECT 91.825 34.740 92.225 35.840 ;
        RECT 93.825 34.740 94.225 35.840 ;
        RECT 95.825 34.740 96.225 35.840 ;
        RECT 97.825 34.740 98.225 35.840 ;
        RECT 99.825 34.740 100.225 35.840 ;
        RECT 101.825 34.740 102.225 35.840 ;
        RECT 103.825 34.740 104.225 35.840 ;
        RECT 105.825 34.740 106.225 35.840 ;
        RECT 107.825 34.740 108.225 35.840 ;
        RECT 109.825 34.740 110.225 35.840 ;
        RECT 111.825 34.740 112.225 35.840 ;
        RECT 113.825 34.740 114.225 35.840 ;
        RECT 115.825 34.740 116.225 35.840 ;
        RECT 117.825 34.740 118.225 35.840 ;
        RECT 119.825 34.740 120.225 35.840 ;
        RECT 121.825 34.740 122.225 35.840 ;
        RECT 123.825 34.740 124.225 35.840 ;
        RECT 125.825 34.740 126.225 35.840 ;
        RECT 127.825 34.740 128.225 35.840 ;
        RECT 129.825 34.740 130.225 35.840 ;
        RECT 131.825 34.740 132.225 35.840 ;
        RECT 133.825 34.740 134.225 35.840 ;
        RECT 135.825 34.740 136.225 35.840 ;
        RECT 137.825 34.740 138.225 35.840 ;
        RECT 139.825 34.740 140.225 35.840 ;
        RECT 141.825 34.740 142.225 35.840 ;
        RECT 143.825 34.740 144.225 35.840 ;
        RECT 145.825 34.740 146.225 35.840 ;
        RECT 147.825 34.740 148.225 35.840 ;
        RECT 149.825 34.740 150.225 35.840 ;
        RECT 151.825 34.740 152.225 35.840 ;
        RECT 153.825 34.740 154.225 35.840 ;
        RECT 87.825 32.890 88.225 33.990 ;
        RECT 89.825 32.890 90.225 33.990 ;
        RECT 91.825 32.890 92.225 33.990 ;
        RECT 93.825 32.890 94.225 33.990 ;
        RECT 95.825 32.890 96.225 33.990 ;
        RECT 97.825 32.890 98.225 33.990 ;
        RECT 99.825 32.890 100.225 33.990 ;
        RECT 101.825 32.890 102.225 33.990 ;
        RECT 103.825 32.890 104.225 33.990 ;
        RECT 105.825 32.890 106.225 33.990 ;
        RECT 107.825 32.890 108.225 33.990 ;
        RECT 109.825 32.890 110.225 33.990 ;
        RECT 111.825 32.890 112.225 33.990 ;
        RECT 113.825 32.890 114.225 33.990 ;
        RECT 115.825 32.890 116.225 33.990 ;
        RECT 117.825 32.890 118.225 33.990 ;
        RECT 119.825 32.890 120.225 33.990 ;
        RECT 121.825 32.890 122.225 33.990 ;
        RECT 123.825 32.890 124.225 33.990 ;
        RECT 125.825 32.890 126.225 33.990 ;
        RECT 127.825 32.890 128.225 33.990 ;
        RECT 129.825 32.890 130.225 33.990 ;
        RECT 131.825 32.890 132.225 33.990 ;
        RECT 133.825 32.890 134.225 33.990 ;
        RECT 135.825 32.890 136.225 33.990 ;
        RECT 137.825 32.890 138.225 33.990 ;
        RECT 139.825 32.890 140.225 33.990 ;
        RECT 141.825 32.890 142.225 33.990 ;
        RECT 143.825 32.890 144.225 33.990 ;
        RECT 145.825 32.890 146.225 33.990 ;
        RECT 147.825 32.890 148.225 33.990 ;
        RECT 149.825 32.890 150.225 33.990 ;
        RECT 151.825 32.890 152.225 33.990 ;
        RECT 153.825 32.890 154.225 33.990 ;
        RECT 87.825 31.040 88.225 32.140 ;
        RECT 89.825 31.040 90.225 32.140 ;
        RECT 91.825 31.040 92.225 32.140 ;
        RECT 93.825 31.040 94.225 32.140 ;
        RECT 95.825 31.040 96.225 32.140 ;
        RECT 97.825 31.040 98.225 32.140 ;
        RECT 99.825 31.040 100.225 32.140 ;
        RECT 101.825 31.040 102.225 32.140 ;
        RECT 103.825 31.040 104.225 32.140 ;
        RECT 105.825 31.040 106.225 32.140 ;
        RECT 107.825 31.040 108.225 32.140 ;
        RECT 109.825 31.040 110.225 32.140 ;
        RECT 111.825 31.040 112.225 32.140 ;
        RECT 113.825 31.040 114.225 32.140 ;
        RECT 115.825 31.040 116.225 32.140 ;
        RECT 117.825 31.040 118.225 32.140 ;
        RECT 119.825 31.040 120.225 32.140 ;
        RECT 121.825 31.040 122.225 32.140 ;
        RECT 123.825 31.040 124.225 32.140 ;
        RECT 125.825 31.040 126.225 32.140 ;
        RECT 127.825 31.040 128.225 32.140 ;
        RECT 129.825 31.040 130.225 32.140 ;
        RECT 131.825 31.040 132.225 32.140 ;
        RECT 133.825 31.040 134.225 32.140 ;
        RECT 135.825 31.040 136.225 32.140 ;
        RECT 137.825 31.040 138.225 32.140 ;
        RECT 139.825 31.040 140.225 32.140 ;
        RECT 141.825 31.040 142.225 32.140 ;
        RECT 143.825 31.040 144.225 32.140 ;
        RECT 145.825 31.040 146.225 32.140 ;
        RECT 147.825 31.040 148.225 32.140 ;
        RECT 149.825 31.040 150.225 32.140 ;
        RECT 151.825 31.040 152.225 32.140 ;
        RECT 153.825 31.040 154.225 32.140 ;
        RECT 87.825 29.190 88.225 30.290 ;
        RECT 89.825 29.190 90.225 30.290 ;
        RECT 91.825 29.190 92.225 30.290 ;
        RECT 93.825 29.190 94.225 30.290 ;
        RECT 95.825 29.190 96.225 30.290 ;
        RECT 97.825 29.190 98.225 30.290 ;
        RECT 99.825 29.190 100.225 30.290 ;
        RECT 101.825 29.190 102.225 30.290 ;
        RECT 103.825 29.190 104.225 30.290 ;
        RECT 105.825 29.190 106.225 30.290 ;
        RECT 107.825 29.190 108.225 30.290 ;
        RECT 109.825 29.190 110.225 30.290 ;
        RECT 111.825 29.190 112.225 30.290 ;
        RECT 113.825 29.190 114.225 30.290 ;
        RECT 115.825 29.190 116.225 30.290 ;
        RECT 117.825 29.190 118.225 30.290 ;
        RECT 119.825 29.190 120.225 30.290 ;
        RECT 121.825 29.190 122.225 30.290 ;
        RECT 123.825 29.190 124.225 30.290 ;
        RECT 125.825 29.190 126.225 30.290 ;
        RECT 127.825 29.190 128.225 30.290 ;
        RECT 129.825 29.190 130.225 30.290 ;
        RECT 131.825 29.190 132.225 30.290 ;
        RECT 133.825 29.190 134.225 30.290 ;
        RECT 135.825 29.190 136.225 30.290 ;
        RECT 137.825 29.190 138.225 30.290 ;
        RECT 139.825 29.190 140.225 30.290 ;
        RECT 141.825 29.190 142.225 30.290 ;
        RECT 143.825 29.190 144.225 30.290 ;
        RECT 145.825 29.190 146.225 30.290 ;
        RECT 147.825 29.190 148.225 30.290 ;
        RECT 149.825 29.190 150.225 30.290 ;
        RECT 151.825 29.190 152.225 30.290 ;
        RECT 153.825 29.190 154.225 30.290 ;
        RECT 87.825 27.340 88.225 28.440 ;
        RECT 89.825 27.340 90.225 28.440 ;
        RECT 91.825 27.340 92.225 28.440 ;
        RECT 93.825 27.340 94.225 28.440 ;
        RECT 95.825 27.340 96.225 28.440 ;
        RECT 97.825 27.340 98.225 28.440 ;
        RECT 99.825 27.340 100.225 28.440 ;
        RECT 101.825 27.340 102.225 28.440 ;
        RECT 103.825 27.340 104.225 28.440 ;
        RECT 105.825 27.340 106.225 28.440 ;
        RECT 107.825 27.340 108.225 28.440 ;
        RECT 109.825 27.340 110.225 28.440 ;
        RECT 111.825 27.340 112.225 28.440 ;
        RECT 113.825 27.340 114.225 28.440 ;
        RECT 115.825 27.340 116.225 28.440 ;
        RECT 117.825 27.340 118.225 28.440 ;
        RECT 119.825 27.340 120.225 28.440 ;
        RECT 121.825 27.340 122.225 28.440 ;
        RECT 123.825 27.340 124.225 28.440 ;
        RECT 125.825 27.340 126.225 28.440 ;
        RECT 127.825 27.340 128.225 28.440 ;
        RECT 129.825 27.340 130.225 28.440 ;
        RECT 131.825 27.340 132.225 28.440 ;
        RECT 133.825 27.340 134.225 28.440 ;
        RECT 135.825 27.340 136.225 28.440 ;
        RECT 137.825 27.340 138.225 28.440 ;
        RECT 139.825 27.340 140.225 28.440 ;
        RECT 141.825 27.340 142.225 28.440 ;
        RECT 143.825 27.340 144.225 28.440 ;
        RECT 145.825 27.340 146.225 28.440 ;
        RECT 147.825 27.340 148.225 28.440 ;
        RECT 149.825 27.340 150.225 28.440 ;
        RECT 151.825 27.340 152.225 28.440 ;
        RECT 153.825 27.340 154.225 28.440 ;
        RECT 74.990 25.840 75.290 26.240 ;
        RECT 85.825 25.840 86.125 26.240 ;
        RECT 87.825 25.490 88.225 26.590 ;
        RECT 89.825 25.490 90.225 26.590 ;
        RECT 91.825 25.490 92.225 26.590 ;
        RECT 93.825 25.490 94.225 26.590 ;
        RECT 95.825 25.490 96.225 26.590 ;
        RECT 97.825 25.490 98.225 26.590 ;
        RECT 99.825 25.490 100.225 26.590 ;
        RECT 101.825 25.490 102.225 26.590 ;
        RECT 103.825 25.490 104.225 26.590 ;
        RECT 105.825 25.490 106.225 26.590 ;
        RECT 107.825 25.490 108.225 26.590 ;
        RECT 109.825 25.490 110.225 26.590 ;
        RECT 111.825 25.490 112.225 26.590 ;
        RECT 113.825 25.490 114.225 26.590 ;
        RECT 115.825 25.490 116.225 26.590 ;
        RECT 117.825 25.490 118.225 26.590 ;
        RECT 119.825 25.490 120.225 26.590 ;
        RECT 121.825 25.490 122.225 26.590 ;
        RECT 123.825 25.490 124.225 26.590 ;
        RECT 125.825 25.490 126.225 26.590 ;
        RECT 127.825 25.490 128.225 26.590 ;
        RECT 129.825 25.490 130.225 26.590 ;
        RECT 131.825 25.490 132.225 26.590 ;
        RECT 133.825 25.490 134.225 26.590 ;
        RECT 135.825 25.490 136.225 26.590 ;
        RECT 137.825 25.490 138.225 26.590 ;
        RECT 139.825 25.490 140.225 26.590 ;
        RECT 141.825 25.490 142.225 26.590 ;
        RECT 143.825 25.490 144.225 26.590 ;
        RECT 145.825 25.490 146.225 26.590 ;
        RECT 147.825 25.490 148.225 26.590 ;
        RECT 149.825 25.490 150.225 26.590 ;
        RECT 151.825 25.490 152.225 26.590 ;
        RECT 153.825 25.490 154.225 26.590 ;
        RECT 6.890 23.640 7.290 24.740 ;
        RECT 8.890 23.640 9.290 24.740 ;
        RECT 10.890 23.640 11.290 24.740 ;
        RECT 12.890 23.640 13.290 24.740 ;
        RECT 14.890 23.640 15.290 24.740 ;
        RECT 16.890 23.640 17.290 24.740 ;
        RECT 18.890 23.640 19.290 24.740 ;
        RECT 20.890 23.640 21.290 24.740 ;
        RECT 22.890 23.640 23.290 24.740 ;
        RECT 24.890 23.640 25.290 24.740 ;
        RECT 26.890 23.640 27.290 24.740 ;
        RECT 28.890 23.640 29.290 24.740 ;
        RECT 30.890 23.640 31.290 24.740 ;
        RECT 32.890 23.640 33.290 24.740 ;
        RECT 34.890 23.640 35.290 24.740 ;
        RECT 36.890 23.640 37.290 24.740 ;
        RECT 38.890 23.640 39.290 24.740 ;
        RECT 40.890 23.640 41.290 24.740 ;
        RECT 42.890 23.640 43.290 24.740 ;
        RECT 44.890 23.640 45.290 24.740 ;
        RECT 46.890 23.640 47.290 24.740 ;
        RECT 48.890 23.640 49.290 24.740 ;
        RECT 50.890 23.640 51.290 24.740 ;
        RECT 52.890 23.640 53.290 24.740 ;
        RECT 54.890 23.640 55.290 24.740 ;
        RECT 56.890 23.640 57.290 24.740 ;
        RECT 58.890 23.640 59.290 24.740 ;
        RECT 60.890 23.640 61.290 24.740 ;
        RECT 62.890 23.640 63.290 24.740 ;
        RECT 64.890 23.640 65.290 24.740 ;
        RECT 66.890 23.640 67.290 24.740 ;
        RECT 68.890 23.640 69.290 24.740 ;
        RECT 70.890 23.640 71.290 24.740 ;
        RECT 72.890 23.640 73.290 24.740 ;
        RECT 87.825 23.640 88.225 24.740 ;
        RECT 89.825 23.640 90.225 24.740 ;
        RECT 91.825 23.640 92.225 24.740 ;
        RECT 93.825 23.640 94.225 24.740 ;
        RECT 95.825 23.640 96.225 24.740 ;
        RECT 97.825 23.640 98.225 24.740 ;
        RECT 99.825 23.640 100.225 24.740 ;
        RECT 101.825 23.640 102.225 24.740 ;
        RECT 103.825 23.640 104.225 24.740 ;
        RECT 105.825 23.640 106.225 24.740 ;
        RECT 107.825 23.640 108.225 24.740 ;
        RECT 109.825 23.640 110.225 24.740 ;
        RECT 111.825 23.640 112.225 24.740 ;
        RECT 113.825 23.640 114.225 24.740 ;
        RECT 115.825 23.640 116.225 24.740 ;
        RECT 117.825 23.640 118.225 24.740 ;
        RECT 119.825 23.640 120.225 24.740 ;
        RECT 121.825 23.640 122.225 24.740 ;
        RECT 123.825 23.640 124.225 24.740 ;
        RECT 125.825 23.640 126.225 24.740 ;
        RECT 127.825 23.640 128.225 24.740 ;
        RECT 129.825 23.640 130.225 24.740 ;
        RECT 131.825 23.640 132.225 24.740 ;
        RECT 133.825 23.640 134.225 24.740 ;
        RECT 135.825 23.640 136.225 24.740 ;
        RECT 137.825 23.640 138.225 24.740 ;
        RECT 139.825 23.640 140.225 24.740 ;
        RECT 141.825 23.640 142.225 24.740 ;
        RECT 143.825 23.640 144.225 24.740 ;
        RECT 145.825 23.640 146.225 24.740 ;
        RECT 147.825 23.640 148.225 24.740 ;
        RECT 149.825 23.640 150.225 24.740 ;
        RECT 151.825 23.640 152.225 24.740 ;
        RECT 153.825 23.640 154.225 24.740 ;
        RECT 6.890 21.790 7.290 22.890 ;
        RECT 8.890 21.790 9.290 22.890 ;
        RECT 10.890 21.790 11.290 22.890 ;
        RECT 12.890 21.790 13.290 22.890 ;
        RECT 14.890 21.790 15.290 22.890 ;
        RECT 16.890 21.790 17.290 22.890 ;
        RECT 18.890 21.790 19.290 22.890 ;
        RECT 20.890 21.790 21.290 22.890 ;
        RECT 22.890 21.790 23.290 22.890 ;
        RECT 24.890 21.790 25.290 22.890 ;
        RECT 26.890 21.790 27.290 22.890 ;
        RECT 28.890 21.790 29.290 22.890 ;
        RECT 30.890 21.790 31.290 22.890 ;
        RECT 32.890 21.790 33.290 22.890 ;
        RECT 34.890 21.790 35.290 22.890 ;
        RECT 36.890 21.790 37.290 22.890 ;
        RECT 38.890 21.790 39.290 22.890 ;
        RECT 40.890 21.790 41.290 22.890 ;
        RECT 42.890 21.790 43.290 22.890 ;
        RECT 44.890 21.790 45.290 22.890 ;
        RECT 46.890 21.790 47.290 22.890 ;
        RECT 48.890 21.790 49.290 22.890 ;
        RECT 50.890 21.790 51.290 22.890 ;
        RECT 52.890 21.790 53.290 22.890 ;
        RECT 54.890 21.790 55.290 22.890 ;
        RECT 56.890 21.790 57.290 22.890 ;
        RECT 58.890 21.790 59.290 22.890 ;
        RECT 60.890 21.790 61.290 22.890 ;
        RECT 62.890 21.790 63.290 22.890 ;
        RECT 64.890 21.790 65.290 22.890 ;
        RECT 66.890 21.790 67.290 22.890 ;
        RECT 68.890 21.790 69.290 22.890 ;
        RECT 70.890 21.790 71.290 22.890 ;
        RECT 72.890 21.790 73.290 22.890 ;
        RECT 87.825 21.790 88.225 22.890 ;
        RECT 89.825 21.790 90.225 22.890 ;
        RECT 91.825 21.790 92.225 22.890 ;
        RECT 93.825 21.790 94.225 22.890 ;
        RECT 95.825 21.790 96.225 22.890 ;
        RECT 97.825 21.790 98.225 22.890 ;
        RECT 99.825 21.790 100.225 22.890 ;
        RECT 101.825 21.790 102.225 22.890 ;
        RECT 103.825 21.790 104.225 22.890 ;
        RECT 105.825 21.790 106.225 22.890 ;
        RECT 107.825 21.790 108.225 22.890 ;
        RECT 109.825 21.790 110.225 22.890 ;
        RECT 111.825 21.790 112.225 22.890 ;
        RECT 113.825 21.790 114.225 22.890 ;
        RECT 115.825 21.790 116.225 22.890 ;
        RECT 117.825 21.790 118.225 22.890 ;
        RECT 119.825 21.790 120.225 22.890 ;
        RECT 121.825 21.790 122.225 22.890 ;
        RECT 123.825 21.790 124.225 22.890 ;
        RECT 125.825 21.790 126.225 22.890 ;
        RECT 127.825 21.790 128.225 22.890 ;
        RECT 129.825 21.790 130.225 22.890 ;
        RECT 131.825 21.790 132.225 22.890 ;
        RECT 133.825 21.790 134.225 22.890 ;
        RECT 135.825 21.790 136.225 22.890 ;
        RECT 137.825 21.790 138.225 22.890 ;
        RECT 139.825 21.790 140.225 22.890 ;
        RECT 141.825 21.790 142.225 22.890 ;
        RECT 143.825 21.790 144.225 22.890 ;
        RECT 145.825 21.790 146.225 22.890 ;
        RECT 147.825 21.790 148.225 22.890 ;
        RECT 149.825 21.790 150.225 22.890 ;
        RECT 151.825 21.790 152.225 22.890 ;
        RECT 153.825 21.790 154.225 22.890 ;
        RECT 6.890 19.940 7.290 21.040 ;
        RECT 8.890 19.940 9.290 21.040 ;
        RECT 10.890 19.940 11.290 21.040 ;
        RECT 12.890 19.940 13.290 21.040 ;
        RECT 14.890 19.940 15.290 21.040 ;
        RECT 16.890 19.940 17.290 21.040 ;
        RECT 18.890 19.940 19.290 21.040 ;
        RECT 20.890 19.940 21.290 21.040 ;
        RECT 22.890 19.940 23.290 21.040 ;
        RECT 24.890 19.940 25.290 21.040 ;
        RECT 26.890 19.940 27.290 21.040 ;
        RECT 28.890 19.940 29.290 21.040 ;
        RECT 30.890 19.940 31.290 21.040 ;
        RECT 32.890 19.940 33.290 21.040 ;
        RECT 34.890 19.940 35.290 21.040 ;
        RECT 36.890 19.940 37.290 21.040 ;
        RECT 38.890 19.940 39.290 21.040 ;
        RECT 40.890 19.940 41.290 21.040 ;
        RECT 42.890 19.940 43.290 21.040 ;
        RECT 44.890 19.940 45.290 21.040 ;
        RECT 46.890 19.940 47.290 21.040 ;
        RECT 48.890 19.940 49.290 21.040 ;
        RECT 50.890 19.940 51.290 21.040 ;
        RECT 52.890 19.940 53.290 21.040 ;
        RECT 54.890 19.940 55.290 21.040 ;
        RECT 56.890 19.940 57.290 21.040 ;
        RECT 58.890 19.940 59.290 21.040 ;
        RECT 60.890 19.940 61.290 21.040 ;
        RECT 62.890 19.940 63.290 21.040 ;
        RECT 64.890 19.940 65.290 21.040 ;
        RECT 66.890 19.940 67.290 21.040 ;
        RECT 68.890 19.940 69.290 21.040 ;
        RECT 70.890 19.940 71.290 21.040 ;
        RECT 72.890 19.940 73.290 21.040 ;
        RECT 87.825 19.940 88.225 21.040 ;
        RECT 89.825 19.940 90.225 21.040 ;
        RECT 91.825 19.940 92.225 21.040 ;
        RECT 93.825 19.940 94.225 21.040 ;
        RECT 95.825 19.940 96.225 21.040 ;
        RECT 97.825 19.940 98.225 21.040 ;
        RECT 99.825 19.940 100.225 21.040 ;
        RECT 101.825 19.940 102.225 21.040 ;
        RECT 103.825 19.940 104.225 21.040 ;
        RECT 105.825 19.940 106.225 21.040 ;
        RECT 107.825 19.940 108.225 21.040 ;
        RECT 109.825 19.940 110.225 21.040 ;
        RECT 111.825 19.940 112.225 21.040 ;
        RECT 113.825 19.940 114.225 21.040 ;
        RECT 115.825 19.940 116.225 21.040 ;
        RECT 117.825 19.940 118.225 21.040 ;
        RECT 119.825 19.940 120.225 21.040 ;
        RECT 121.825 19.940 122.225 21.040 ;
        RECT 123.825 19.940 124.225 21.040 ;
        RECT 125.825 19.940 126.225 21.040 ;
        RECT 127.825 19.940 128.225 21.040 ;
        RECT 129.825 19.940 130.225 21.040 ;
        RECT 131.825 19.940 132.225 21.040 ;
        RECT 133.825 19.940 134.225 21.040 ;
        RECT 135.825 19.940 136.225 21.040 ;
        RECT 137.825 19.940 138.225 21.040 ;
        RECT 139.825 19.940 140.225 21.040 ;
        RECT 141.825 19.940 142.225 21.040 ;
        RECT 143.825 19.940 144.225 21.040 ;
        RECT 145.825 19.940 146.225 21.040 ;
        RECT 147.825 19.940 148.225 21.040 ;
        RECT 149.825 19.940 150.225 21.040 ;
        RECT 151.825 19.940 152.225 21.040 ;
        RECT 153.825 19.940 154.225 21.040 ;
        RECT 6.890 18.090 7.290 19.190 ;
        RECT 8.890 18.090 9.290 19.190 ;
        RECT 10.890 18.090 11.290 19.190 ;
        RECT 12.890 18.090 13.290 19.190 ;
        RECT 14.890 18.090 15.290 19.190 ;
        RECT 16.890 18.090 17.290 19.190 ;
        RECT 18.890 18.090 19.290 19.190 ;
        RECT 20.890 18.090 21.290 19.190 ;
        RECT 22.890 18.090 23.290 19.190 ;
        RECT 24.890 18.090 25.290 19.190 ;
        RECT 26.890 18.090 27.290 19.190 ;
        RECT 28.890 18.090 29.290 19.190 ;
        RECT 30.890 18.090 31.290 19.190 ;
        RECT 32.890 18.090 33.290 19.190 ;
        RECT 34.890 18.090 35.290 19.190 ;
        RECT 36.890 18.090 37.290 19.190 ;
        RECT 38.890 18.090 39.290 19.190 ;
        RECT 40.890 18.090 41.290 19.190 ;
        RECT 42.890 18.090 43.290 19.190 ;
        RECT 44.890 18.090 45.290 19.190 ;
        RECT 46.890 18.090 47.290 19.190 ;
        RECT 48.890 18.090 49.290 19.190 ;
        RECT 50.890 18.090 51.290 19.190 ;
        RECT 52.890 18.090 53.290 19.190 ;
        RECT 54.890 18.090 55.290 19.190 ;
        RECT 56.890 18.090 57.290 19.190 ;
        RECT 58.890 18.090 59.290 19.190 ;
        RECT 60.890 18.090 61.290 19.190 ;
        RECT 62.890 18.090 63.290 19.190 ;
        RECT 64.890 18.090 65.290 19.190 ;
        RECT 66.890 18.090 67.290 19.190 ;
        RECT 68.890 18.090 69.290 19.190 ;
        RECT 70.890 18.090 71.290 19.190 ;
        RECT 72.890 18.090 73.290 19.190 ;
        RECT 87.825 18.090 88.225 19.190 ;
        RECT 89.825 18.090 90.225 19.190 ;
        RECT 91.825 18.090 92.225 19.190 ;
        RECT 93.825 18.090 94.225 19.190 ;
        RECT 95.825 18.090 96.225 19.190 ;
        RECT 97.825 18.090 98.225 19.190 ;
        RECT 99.825 18.090 100.225 19.190 ;
        RECT 101.825 18.090 102.225 19.190 ;
        RECT 103.825 18.090 104.225 19.190 ;
        RECT 105.825 18.090 106.225 19.190 ;
        RECT 107.825 18.090 108.225 19.190 ;
        RECT 109.825 18.090 110.225 19.190 ;
        RECT 111.825 18.090 112.225 19.190 ;
        RECT 113.825 18.090 114.225 19.190 ;
        RECT 115.825 18.090 116.225 19.190 ;
        RECT 117.825 18.090 118.225 19.190 ;
        RECT 119.825 18.090 120.225 19.190 ;
        RECT 121.825 18.090 122.225 19.190 ;
        RECT 123.825 18.090 124.225 19.190 ;
        RECT 125.825 18.090 126.225 19.190 ;
        RECT 127.825 18.090 128.225 19.190 ;
        RECT 129.825 18.090 130.225 19.190 ;
        RECT 131.825 18.090 132.225 19.190 ;
        RECT 133.825 18.090 134.225 19.190 ;
        RECT 135.825 18.090 136.225 19.190 ;
        RECT 137.825 18.090 138.225 19.190 ;
        RECT 139.825 18.090 140.225 19.190 ;
        RECT 141.825 18.090 142.225 19.190 ;
        RECT 143.825 18.090 144.225 19.190 ;
        RECT 145.825 18.090 146.225 19.190 ;
        RECT 147.825 18.090 148.225 19.190 ;
        RECT 149.825 18.090 150.225 19.190 ;
        RECT 151.825 18.090 152.225 19.190 ;
        RECT 153.825 18.090 154.225 19.190 ;
        RECT 6.890 16.240 7.290 17.340 ;
        RECT 8.890 16.240 9.290 17.340 ;
        RECT 10.890 16.240 11.290 17.340 ;
        RECT 12.890 16.240 13.290 17.340 ;
        RECT 14.890 16.240 15.290 17.340 ;
        RECT 16.890 16.240 17.290 17.340 ;
        RECT 18.890 16.240 19.290 17.340 ;
        RECT 20.890 16.240 21.290 17.340 ;
        RECT 22.890 16.240 23.290 17.340 ;
        RECT 24.890 16.240 25.290 17.340 ;
        RECT 26.890 16.240 27.290 17.340 ;
        RECT 28.890 16.240 29.290 17.340 ;
        RECT 30.890 16.240 31.290 17.340 ;
        RECT 32.890 16.240 33.290 17.340 ;
        RECT 34.890 16.240 35.290 17.340 ;
        RECT 36.890 16.240 37.290 17.340 ;
        RECT 38.890 16.240 39.290 17.340 ;
        RECT 40.890 16.240 41.290 17.340 ;
        RECT 42.890 16.240 43.290 17.340 ;
        RECT 44.890 16.240 45.290 17.340 ;
        RECT 46.890 16.240 47.290 17.340 ;
        RECT 48.890 16.240 49.290 17.340 ;
        RECT 50.890 16.240 51.290 17.340 ;
        RECT 52.890 16.240 53.290 17.340 ;
        RECT 54.890 16.240 55.290 17.340 ;
        RECT 56.890 16.240 57.290 17.340 ;
        RECT 58.890 16.240 59.290 17.340 ;
        RECT 60.890 16.240 61.290 17.340 ;
        RECT 62.890 16.240 63.290 17.340 ;
        RECT 64.890 16.240 65.290 17.340 ;
        RECT 66.890 16.240 67.290 17.340 ;
        RECT 68.890 16.240 69.290 17.340 ;
        RECT 70.890 16.240 71.290 17.340 ;
        RECT 72.890 16.240 73.290 17.340 ;
        RECT 87.825 16.240 88.225 17.340 ;
        RECT 89.825 16.240 90.225 17.340 ;
        RECT 91.825 16.240 92.225 17.340 ;
        RECT 93.825 16.240 94.225 17.340 ;
        RECT 95.825 16.240 96.225 17.340 ;
        RECT 97.825 16.240 98.225 17.340 ;
        RECT 99.825 16.240 100.225 17.340 ;
        RECT 101.825 16.240 102.225 17.340 ;
        RECT 103.825 16.240 104.225 17.340 ;
        RECT 105.825 16.240 106.225 17.340 ;
        RECT 107.825 16.240 108.225 17.340 ;
        RECT 109.825 16.240 110.225 17.340 ;
        RECT 111.825 16.240 112.225 17.340 ;
        RECT 113.825 16.240 114.225 17.340 ;
        RECT 115.825 16.240 116.225 17.340 ;
        RECT 117.825 16.240 118.225 17.340 ;
        RECT 119.825 16.240 120.225 17.340 ;
        RECT 121.825 16.240 122.225 17.340 ;
        RECT 123.825 16.240 124.225 17.340 ;
        RECT 125.825 16.240 126.225 17.340 ;
        RECT 127.825 16.240 128.225 17.340 ;
        RECT 129.825 16.240 130.225 17.340 ;
        RECT 131.825 16.240 132.225 17.340 ;
        RECT 133.825 16.240 134.225 17.340 ;
        RECT 135.825 16.240 136.225 17.340 ;
        RECT 137.825 16.240 138.225 17.340 ;
        RECT 139.825 16.240 140.225 17.340 ;
        RECT 141.825 16.240 142.225 17.340 ;
        RECT 143.825 16.240 144.225 17.340 ;
        RECT 145.825 16.240 146.225 17.340 ;
        RECT 147.825 16.240 148.225 17.340 ;
        RECT 149.825 16.240 150.225 17.340 ;
        RECT 151.825 16.240 152.225 17.340 ;
        RECT 153.825 16.240 154.225 17.340 ;
        RECT 6.890 14.390 7.290 15.490 ;
        RECT 8.890 14.390 9.290 15.490 ;
        RECT 10.890 14.390 11.290 15.490 ;
        RECT 12.890 14.390 13.290 15.490 ;
        RECT 14.890 14.390 15.290 15.490 ;
        RECT 16.890 14.390 17.290 15.490 ;
        RECT 18.890 14.390 19.290 15.490 ;
        RECT 20.890 14.390 21.290 15.490 ;
        RECT 22.890 14.390 23.290 15.490 ;
        RECT 24.890 14.390 25.290 15.490 ;
        RECT 26.890 14.390 27.290 15.490 ;
        RECT 28.890 14.390 29.290 15.490 ;
        RECT 30.890 14.390 31.290 15.490 ;
        RECT 32.890 14.390 33.290 15.490 ;
        RECT 34.890 14.390 35.290 15.490 ;
        RECT 36.890 14.390 37.290 15.490 ;
        RECT 38.890 14.390 39.290 15.490 ;
        RECT 40.890 14.390 41.290 15.490 ;
        RECT 42.890 14.390 43.290 15.490 ;
        RECT 44.890 14.390 45.290 15.490 ;
        RECT 46.890 14.390 47.290 15.490 ;
        RECT 48.890 14.390 49.290 15.490 ;
        RECT 50.890 14.390 51.290 15.490 ;
        RECT 52.890 14.390 53.290 15.490 ;
        RECT 54.890 14.390 55.290 15.490 ;
        RECT 56.890 14.390 57.290 15.490 ;
        RECT 58.890 14.390 59.290 15.490 ;
        RECT 60.890 14.390 61.290 15.490 ;
        RECT 62.890 14.390 63.290 15.490 ;
        RECT 64.890 14.390 65.290 15.490 ;
        RECT 66.890 14.390 67.290 15.490 ;
        RECT 68.890 14.390 69.290 15.490 ;
        RECT 70.890 14.390 71.290 15.490 ;
        RECT 72.890 14.390 73.290 15.490 ;
        RECT 87.825 14.390 88.225 15.490 ;
        RECT 89.825 14.390 90.225 15.490 ;
        RECT 91.825 14.390 92.225 15.490 ;
        RECT 93.825 14.390 94.225 15.490 ;
        RECT 95.825 14.390 96.225 15.490 ;
        RECT 97.825 14.390 98.225 15.490 ;
        RECT 99.825 14.390 100.225 15.490 ;
        RECT 101.825 14.390 102.225 15.490 ;
        RECT 103.825 14.390 104.225 15.490 ;
        RECT 105.825 14.390 106.225 15.490 ;
        RECT 107.825 14.390 108.225 15.490 ;
        RECT 109.825 14.390 110.225 15.490 ;
        RECT 111.825 14.390 112.225 15.490 ;
        RECT 113.825 14.390 114.225 15.490 ;
        RECT 115.825 14.390 116.225 15.490 ;
        RECT 117.825 14.390 118.225 15.490 ;
        RECT 119.825 14.390 120.225 15.490 ;
        RECT 121.825 14.390 122.225 15.490 ;
        RECT 123.825 14.390 124.225 15.490 ;
        RECT 125.825 14.390 126.225 15.490 ;
        RECT 127.825 14.390 128.225 15.490 ;
        RECT 129.825 14.390 130.225 15.490 ;
        RECT 131.825 14.390 132.225 15.490 ;
        RECT 133.825 14.390 134.225 15.490 ;
        RECT 135.825 14.390 136.225 15.490 ;
        RECT 137.825 14.390 138.225 15.490 ;
        RECT 139.825 14.390 140.225 15.490 ;
        RECT 141.825 14.390 142.225 15.490 ;
        RECT 143.825 14.390 144.225 15.490 ;
        RECT 145.825 14.390 146.225 15.490 ;
        RECT 147.825 14.390 148.225 15.490 ;
        RECT 149.825 14.390 150.225 15.490 ;
        RECT 151.825 14.390 152.225 15.490 ;
        RECT 153.825 14.390 154.225 15.490 ;
        RECT 6.890 12.540 7.290 13.640 ;
        RECT 8.890 12.540 9.290 13.640 ;
        RECT 10.890 12.540 11.290 13.640 ;
        RECT 12.890 12.540 13.290 13.640 ;
        RECT 14.890 12.540 15.290 13.640 ;
        RECT 16.890 12.540 17.290 13.640 ;
        RECT 18.890 12.540 19.290 13.640 ;
        RECT 20.890 12.540 21.290 13.640 ;
        RECT 22.890 12.540 23.290 13.640 ;
        RECT 24.890 12.540 25.290 13.640 ;
        RECT 26.890 12.540 27.290 13.640 ;
        RECT 28.890 12.540 29.290 13.640 ;
        RECT 30.890 12.540 31.290 13.640 ;
        RECT 32.890 12.540 33.290 13.640 ;
        RECT 34.890 12.540 35.290 13.640 ;
        RECT 36.890 12.540 37.290 13.640 ;
        RECT 38.890 12.540 39.290 13.640 ;
        RECT 40.890 12.540 41.290 13.640 ;
        RECT 42.890 12.540 43.290 13.640 ;
        RECT 44.890 12.540 45.290 13.640 ;
        RECT 46.890 12.540 47.290 13.640 ;
        RECT 48.890 12.540 49.290 13.640 ;
        RECT 50.890 12.540 51.290 13.640 ;
        RECT 52.890 12.540 53.290 13.640 ;
        RECT 54.890 12.540 55.290 13.640 ;
        RECT 56.890 12.540 57.290 13.640 ;
        RECT 58.890 12.540 59.290 13.640 ;
        RECT 60.890 12.540 61.290 13.640 ;
        RECT 62.890 12.540 63.290 13.640 ;
        RECT 64.890 12.540 65.290 13.640 ;
        RECT 66.890 12.540 67.290 13.640 ;
        RECT 68.890 12.540 69.290 13.640 ;
        RECT 70.890 12.540 71.290 13.640 ;
        RECT 72.890 12.540 73.290 13.640 ;
        RECT 87.825 12.540 88.225 13.640 ;
        RECT 89.825 12.540 90.225 13.640 ;
        RECT 91.825 12.540 92.225 13.640 ;
        RECT 93.825 12.540 94.225 13.640 ;
        RECT 95.825 12.540 96.225 13.640 ;
        RECT 97.825 12.540 98.225 13.640 ;
        RECT 99.825 12.540 100.225 13.640 ;
        RECT 101.825 12.540 102.225 13.640 ;
        RECT 103.825 12.540 104.225 13.640 ;
        RECT 105.825 12.540 106.225 13.640 ;
        RECT 107.825 12.540 108.225 13.640 ;
        RECT 109.825 12.540 110.225 13.640 ;
        RECT 111.825 12.540 112.225 13.640 ;
        RECT 113.825 12.540 114.225 13.640 ;
        RECT 115.825 12.540 116.225 13.640 ;
        RECT 117.825 12.540 118.225 13.640 ;
        RECT 119.825 12.540 120.225 13.640 ;
        RECT 121.825 12.540 122.225 13.640 ;
        RECT 123.825 12.540 124.225 13.640 ;
        RECT 125.825 12.540 126.225 13.640 ;
        RECT 127.825 12.540 128.225 13.640 ;
        RECT 129.825 12.540 130.225 13.640 ;
        RECT 131.825 12.540 132.225 13.640 ;
        RECT 133.825 12.540 134.225 13.640 ;
        RECT 135.825 12.540 136.225 13.640 ;
        RECT 137.825 12.540 138.225 13.640 ;
        RECT 139.825 12.540 140.225 13.640 ;
        RECT 141.825 12.540 142.225 13.640 ;
        RECT 143.825 12.540 144.225 13.640 ;
        RECT 145.825 12.540 146.225 13.640 ;
        RECT 147.825 12.540 148.225 13.640 ;
        RECT 149.825 12.540 150.225 13.640 ;
        RECT 151.825 12.540 152.225 13.640 ;
        RECT 153.825 12.540 154.225 13.640 ;
        RECT 6.890 10.690 7.290 11.790 ;
        RECT 8.890 10.690 9.290 11.790 ;
        RECT 10.890 10.690 11.290 11.790 ;
        RECT 12.890 10.690 13.290 11.790 ;
        RECT 14.890 10.690 15.290 11.790 ;
        RECT 16.890 10.690 17.290 11.790 ;
        RECT 18.890 10.690 19.290 11.790 ;
        RECT 20.890 10.690 21.290 11.790 ;
        RECT 22.890 10.690 23.290 11.790 ;
        RECT 24.890 10.690 25.290 11.790 ;
        RECT 26.890 10.690 27.290 11.790 ;
        RECT 28.890 10.690 29.290 11.790 ;
        RECT 30.890 10.690 31.290 11.790 ;
        RECT 32.890 10.690 33.290 11.790 ;
        RECT 34.890 10.690 35.290 11.790 ;
        RECT 36.890 10.690 37.290 11.790 ;
        RECT 38.890 10.690 39.290 11.790 ;
        RECT 40.890 10.690 41.290 11.790 ;
        RECT 42.890 10.690 43.290 11.790 ;
        RECT 44.890 10.690 45.290 11.790 ;
        RECT 46.890 10.690 47.290 11.790 ;
        RECT 48.890 10.690 49.290 11.790 ;
        RECT 50.890 10.690 51.290 11.790 ;
        RECT 52.890 10.690 53.290 11.790 ;
        RECT 54.890 10.690 55.290 11.790 ;
        RECT 56.890 10.690 57.290 11.790 ;
        RECT 58.890 10.690 59.290 11.790 ;
        RECT 60.890 10.690 61.290 11.790 ;
        RECT 62.890 10.690 63.290 11.790 ;
        RECT 64.890 10.690 65.290 11.790 ;
        RECT 66.890 10.690 67.290 11.790 ;
        RECT 68.890 10.690 69.290 11.790 ;
        RECT 70.890 10.690 71.290 11.790 ;
        RECT 72.890 10.690 73.290 11.790 ;
        RECT 87.825 10.690 88.225 11.790 ;
        RECT 89.825 10.690 90.225 11.790 ;
        RECT 91.825 10.690 92.225 11.790 ;
        RECT 93.825 10.690 94.225 11.790 ;
        RECT 95.825 10.690 96.225 11.790 ;
        RECT 97.825 10.690 98.225 11.790 ;
        RECT 99.825 10.690 100.225 11.790 ;
        RECT 101.825 10.690 102.225 11.790 ;
        RECT 103.825 10.690 104.225 11.790 ;
        RECT 105.825 10.690 106.225 11.790 ;
        RECT 107.825 10.690 108.225 11.790 ;
        RECT 109.825 10.690 110.225 11.790 ;
        RECT 111.825 10.690 112.225 11.790 ;
        RECT 113.825 10.690 114.225 11.790 ;
        RECT 115.825 10.690 116.225 11.790 ;
        RECT 117.825 10.690 118.225 11.790 ;
        RECT 119.825 10.690 120.225 11.790 ;
        RECT 121.825 10.690 122.225 11.790 ;
        RECT 123.825 10.690 124.225 11.790 ;
        RECT 125.825 10.690 126.225 11.790 ;
        RECT 127.825 10.690 128.225 11.790 ;
        RECT 129.825 10.690 130.225 11.790 ;
        RECT 131.825 10.690 132.225 11.790 ;
        RECT 133.825 10.690 134.225 11.790 ;
        RECT 135.825 10.690 136.225 11.790 ;
        RECT 137.825 10.690 138.225 11.790 ;
        RECT 139.825 10.690 140.225 11.790 ;
        RECT 141.825 10.690 142.225 11.790 ;
        RECT 143.825 10.690 144.225 11.790 ;
        RECT 145.825 10.690 146.225 11.790 ;
        RECT 147.825 10.690 148.225 11.790 ;
        RECT 149.825 10.690 150.225 11.790 ;
        RECT 151.825 10.690 152.225 11.790 ;
        RECT 153.825 10.690 154.225 11.790 ;
        RECT 6.890 8.840 7.290 9.940 ;
        RECT 8.890 8.840 9.290 9.940 ;
        RECT 10.890 8.840 11.290 9.940 ;
        RECT 12.890 8.840 13.290 9.940 ;
        RECT 14.890 8.840 15.290 9.940 ;
        RECT 16.890 8.840 17.290 9.940 ;
        RECT 18.890 8.840 19.290 9.940 ;
        RECT 20.890 8.840 21.290 9.940 ;
        RECT 22.890 8.840 23.290 9.940 ;
        RECT 24.890 8.840 25.290 9.940 ;
        RECT 26.890 8.840 27.290 9.940 ;
        RECT 28.890 8.840 29.290 9.940 ;
        RECT 30.890 8.840 31.290 9.940 ;
        RECT 32.890 8.840 33.290 9.940 ;
        RECT 34.890 8.840 35.290 9.940 ;
        RECT 36.890 8.840 37.290 9.940 ;
        RECT 38.890 8.840 39.290 9.940 ;
        RECT 40.890 8.840 41.290 9.940 ;
        RECT 42.890 8.840 43.290 9.940 ;
        RECT 44.890 8.840 45.290 9.940 ;
        RECT 46.890 8.840 47.290 9.940 ;
        RECT 48.890 8.840 49.290 9.940 ;
        RECT 50.890 8.840 51.290 9.940 ;
        RECT 52.890 8.840 53.290 9.940 ;
        RECT 54.890 8.840 55.290 9.940 ;
        RECT 56.890 8.840 57.290 9.940 ;
        RECT 58.890 8.840 59.290 9.940 ;
        RECT 60.890 8.840 61.290 9.940 ;
        RECT 62.890 8.840 63.290 9.940 ;
        RECT 64.890 8.840 65.290 9.940 ;
        RECT 66.890 8.840 67.290 9.940 ;
        RECT 68.890 8.840 69.290 9.940 ;
        RECT 70.890 8.840 71.290 9.940 ;
        RECT 72.890 8.840 73.290 9.940 ;
        RECT 87.825 8.840 88.225 9.940 ;
        RECT 89.825 8.840 90.225 9.940 ;
        RECT 91.825 8.840 92.225 9.940 ;
        RECT 93.825 8.840 94.225 9.940 ;
        RECT 95.825 8.840 96.225 9.940 ;
        RECT 97.825 8.840 98.225 9.940 ;
        RECT 99.825 8.840 100.225 9.940 ;
        RECT 101.825 8.840 102.225 9.940 ;
        RECT 103.825 8.840 104.225 9.940 ;
        RECT 105.825 8.840 106.225 9.940 ;
        RECT 107.825 8.840 108.225 9.940 ;
        RECT 109.825 8.840 110.225 9.940 ;
        RECT 111.825 8.840 112.225 9.940 ;
        RECT 113.825 8.840 114.225 9.940 ;
        RECT 115.825 8.840 116.225 9.940 ;
        RECT 117.825 8.840 118.225 9.940 ;
        RECT 119.825 8.840 120.225 9.940 ;
        RECT 121.825 8.840 122.225 9.940 ;
        RECT 123.825 8.840 124.225 9.940 ;
        RECT 125.825 8.840 126.225 9.940 ;
        RECT 127.825 8.840 128.225 9.940 ;
        RECT 129.825 8.840 130.225 9.940 ;
        RECT 131.825 8.840 132.225 9.940 ;
        RECT 133.825 8.840 134.225 9.940 ;
        RECT 135.825 8.840 136.225 9.940 ;
        RECT 137.825 8.840 138.225 9.940 ;
        RECT 139.825 8.840 140.225 9.940 ;
        RECT 141.825 8.840 142.225 9.940 ;
        RECT 143.825 8.840 144.225 9.940 ;
        RECT 145.825 8.840 146.225 9.940 ;
        RECT 147.825 8.840 148.225 9.940 ;
        RECT 149.825 8.840 150.225 9.940 ;
        RECT 151.825 8.840 152.225 9.940 ;
        RECT 153.825 8.840 154.225 9.940 ;
        RECT 6.890 6.990 7.290 8.090 ;
        RECT 8.890 6.990 9.290 8.090 ;
        RECT 10.890 6.990 11.290 8.090 ;
        RECT 12.890 6.990 13.290 8.090 ;
        RECT 14.890 6.990 15.290 8.090 ;
        RECT 16.890 6.990 17.290 8.090 ;
        RECT 18.890 6.990 19.290 8.090 ;
        RECT 20.890 6.990 21.290 8.090 ;
        RECT 22.890 6.990 23.290 8.090 ;
        RECT 24.890 6.990 25.290 8.090 ;
        RECT 26.890 6.990 27.290 8.090 ;
        RECT 28.890 6.990 29.290 8.090 ;
        RECT 30.890 6.990 31.290 8.090 ;
        RECT 32.890 6.990 33.290 8.090 ;
        RECT 34.890 6.990 35.290 8.090 ;
        RECT 36.890 6.990 37.290 8.090 ;
        RECT 38.890 6.990 39.290 8.090 ;
        RECT 40.890 6.990 41.290 8.090 ;
        RECT 42.890 6.990 43.290 8.090 ;
        RECT 44.890 6.990 45.290 8.090 ;
        RECT 46.890 6.990 47.290 8.090 ;
        RECT 48.890 6.990 49.290 8.090 ;
        RECT 50.890 6.990 51.290 8.090 ;
        RECT 52.890 6.990 53.290 8.090 ;
        RECT 54.890 6.990 55.290 8.090 ;
        RECT 56.890 6.990 57.290 8.090 ;
        RECT 58.890 6.990 59.290 8.090 ;
        RECT 60.890 6.990 61.290 8.090 ;
        RECT 62.890 6.990 63.290 8.090 ;
        RECT 64.890 6.990 65.290 8.090 ;
        RECT 66.890 6.990 67.290 8.090 ;
        RECT 68.890 6.990 69.290 8.090 ;
        RECT 70.890 6.990 71.290 8.090 ;
        RECT 72.890 6.990 73.290 8.090 ;
        RECT 87.825 6.990 88.225 8.090 ;
        RECT 89.825 6.990 90.225 8.090 ;
        RECT 91.825 6.990 92.225 8.090 ;
        RECT 93.825 6.990 94.225 8.090 ;
        RECT 95.825 6.990 96.225 8.090 ;
        RECT 97.825 6.990 98.225 8.090 ;
        RECT 99.825 6.990 100.225 8.090 ;
        RECT 101.825 6.990 102.225 8.090 ;
        RECT 103.825 6.990 104.225 8.090 ;
        RECT 105.825 6.990 106.225 8.090 ;
        RECT 107.825 6.990 108.225 8.090 ;
        RECT 109.825 6.990 110.225 8.090 ;
        RECT 111.825 6.990 112.225 8.090 ;
        RECT 113.825 6.990 114.225 8.090 ;
        RECT 115.825 6.990 116.225 8.090 ;
        RECT 117.825 6.990 118.225 8.090 ;
        RECT 119.825 6.990 120.225 8.090 ;
        RECT 121.825 6.990 122.225 8.090 ;
        RECT 123.825 6.990 124.225 8.090 ;
        RECT 125.825 6.990 126.225 8.090 ;
        RECT 127.825 6.990 128.225 8.090 ;
        RECT 129.825 6.990 130.225 8.090 ;
        RECT 131.825 6.990 132.225 8.090 ;
        RECT 133.825 6.990 134.225 8.090 ;
        RECT 135.825 6.990 136.225 8.090 ;
        RECT 137.825 6.990 138.225 8.090 ;
        RECT 139.825 6.990 140.225 8.090 ;
        RECT 141.825 6.990 142.225 8.090 ;
        RECT 143.825 6.990 144.225 8.090 ;
        RECT 145.825 6.990 146.225 8.090 ;
        RECT 147.825 6.990 148.225 8.090 ;
        RECT 149.825 6.990 150.225 8.090 ;
        RECT 151.825 6.990 152.225 8.090 ;
        RECT 153.825 6.990 154.225 8.090 ;
        RECT 6.890 5.140 7.290 6.240 ;
        RECT 8.890 5.140 9.290 6.240 ;
        RECT 10.890 5.140 11.290 6.240 ;
        RECT 12.890 5.140 13.290 6.240 ;
        RECT 14.890 5.140 15.290 6.240 ;
        RECT 16.890 5.140 17.290 6.240 ;
        RECT 18.890 5.140 19.290 6.240 ;
        RECT 20.890 5.140 21.290 6.240 ;
        RECT 22.890 5.140 23.290 6.240 ;
        RECT 24.890 5.140 25.290 6.240 ;
        RECT 26.890 5.140 27.290 6.240 ;
        RECT 28.890 5.140 29.290 6.240 ;
        RECT 30.890 5.140 31.290 6.240 ;
        RECT 32.890 5.140 33.290 6.240 ;
        RECT 34.890 5.140 35.290 6.240 ;
        RECT 36.890 5.140 37.290 6.240 ;
        RECT 38.890 5.140 39.290 6.240 ;
        RECT 40.890 5.140 41.290 6.240 ;
        RECT 42.890 5.140 43.290 6.240 ;
        RECT 44.890 5.140 45.290 6.240 ;
        RECT 46.890 5.140 47.290 6.240 ;
        RECT 48.890 5.140 49.290 6.240 ;
        RECT 50.890 5.140 51.290 6.240 ;
        RECT 52.890 5.140 53.290 6.240 ;
        RECT 54.890 5.140 55.290 6.240 ;
        RECT 56.890 5.140 57.290 6.240 ;
        RECT 58.890 5.140 59.290 6.240 ;
        RECT 60.890 5.140 61.290 6.240 ;
        RECT 62.890 5.140 63.290 6.240 ;
        RECT 64.890 5.140 65.290 6.240 ;
        RECT 66.890 5.140 67.290 6.240 ;
        RECT 68.890 5.140 69.290 6.240 ;
        RECT 70.890 5.140 71.290 6.240 ;
        RECT 72.890 5.140 73.290 6.240 ;
        RECT 87.825 5.140 88.225 6.240 ;
        RECT 89.825 5.140 90.225 6.240 ;
        RECT 91.825 5.140 92.225 6.240 ;
        RECT 93.825 5.140 94.225 6.240 ;
        RECT 95.825 5.140 96.225 6.240 ;
        RECT 97.825 5.140 98.225 6.240 ;
        RECT 99.825 5.140 100.225 6.240 ;
        RECT 101.825 5.140 102.225 6.240 ;
        RECT 103.825 5.140 104.225 6.240 ;
        RECT 105.825 5.140 106.225 6.240 ;
        RECT 107.825 5.140 108.225 6.240 ;
        RECT 109.825 5.140 110.225 6.240 ;
        RECT 111.825 5.140 112.225 6.240 ;
        RECT 113.825 5.140 114.225 6.240 ;
        RECT 115.825 5.140 116.225 6.240 ;
        RECT 117.825 5.140 118.225 6.240 ;
        RECT 119.825 5.140 120.225 6.240 ;
        RECT 121.825 5.140 122.225 6.240 ;
        RECT 123.825 5.140 124.225 6.240 ;
        RECT 125.825 5.140 126.225 6.240 ;
        RECT 127.825 5.140 128.225 6.240 ;
        RECT 129.825 5.140 130.225 6.240 ;
        RECT 131.825 5.140 132.225 6.240 ;
        RECT 133.825 5.140 134.225 6.240 ;
        RECT 135.825 5.140 136.225 6.240 ;
        RECT 137.825 5.140 138.225 6.240 ;
        RECT 139.825 5.140 140.225 6.240 ;
        RECT 141.825 5.140 142.225 6.240 ;
        RECT 143.825 5.140 144.225 6.240 ;
        RECT 145.825 5.140 146.225 6.240 ;
        RECT 147.825 5.140 148.225 6.240 ;
        RECT 149.825 5.140 150.225 6.240 ;
        RECT 151.825 5.140 152.225 6.240 ;
        RECT 153.825 5.140 154.225 6.240 ;
      LAYER met3 ;
        RECT 3.900 224.100 4.400 224.150 ;
        RECT 7.550 224.100 8.050 224.150 ;
        RECT 11.250 224.100 11.750 224.150 ;
        RECT 14.900 224.100 15.400 224.150 ;
        RECT 18.600 224.100 19.100 224.150 ;
        RECT 22.300 224.100 22.800 224.150 ;
        RECT 25.950 224.100 26.450 224.150 ;
        RECT 29.650 224.100 30.150 224.150 ;
        RECT 33.350 224.100 33.850 224.150 ;
        RECT 37.000 224.100 37.500 224.150 ;
        RECT 40.700 224.100 41.200 224.150 ;
        RECT 44.400 224.100 44.900 224.150 ;
        RECT 48.050 224.100 48.550 224.150 ;
        RECT 51.700 224.100 52.200 224.150 ;
        RECT 55.400 224.100 55.900 224.150 ;
        RECT 59.100 224.100 59.600 224.150 ;
        RECT 3.900 223.800 159.650 224.100 ;
        RECT 3.900 223.750 4.400 223.800 ;
        RECT 7.550 223.750 8.050 223.800 ;
        RECT 11.250 223.750 11.750 223.800 ;
        RECT 14.900 223.750 15.400 223.800 ;
        RECT 18.600 223.750 19.100 223.800 ;
        RECT 22.300 223.750 22.800 223.800 ;
        RECT 25.950 223.750 26.450 223.800 ;
        RECT 29.650 223.750 30.150 223.800 ;
        RECT 33.350 223.750 33.850 223.800 ;
        RECT 37.000 223.750 37.500 223.800 ;
        RECT 40.700 223.750 41.200 223.800 ;
        RECT 44.400 223.750 44.900 223.800 ;
        RECT 48.050 223.750 48.550 223.800 ;
        RECT 51.700 223.750 52.200 223.800 ;
        RECT 55.400 223.750 55.900 223.800 ;
        RECT 59.100 223.750 59.600 223.800 ;
        RECT 159.150 223.700 159.650 223.800 ;
        RECT 14.800 223.400 15.200 223.450 ;
        RECT 66.400 223.400 66.900 223.500 ;
        RECT 14.800 223.100 66.900 223.400 ;
        RECT 134.400 223.400 134.800 223.425 ;
        RECT 140.020 223.400 140.520 223.500 ;
        RECT 134.400 223.100 140.520 223.400 ;
        RECT 134.400 223.075 134.800 223.100 ;
        RECT 70.100 222.800 70.600 222.900 ;
        RECT 26.760 222.500 70.600 222.800 ;
        RECT 143.700 222.800 144.200 222.900 ;
        RECT 146.350 222.800 146.750 222.875 ;
        RECT 143.700 222.500 146.750 222.800 ;
        RECT 26.760 222.450 27.160 222.500 ;
        RECT 73.750 222.200 74.250 222.300 ;
        RECT 38.720 221.900 74.250 222.200 ;
        RECT 122.450 222.200 122.850 222.300 ;
        RECT 147.380 222.200 147.880 222.300 ;
        RECT 122.450 221.900 147.880 222.200 ;
        RECT 38.720 221.850 39.120 221.900 ;
        RECT 77.500 221.600 78.000 221.700 ;
        RECT 50.680 221.300 78.000 221.600 ;
        RECT 98.550 221.600 98.950 221.625 ;
        RECT 151.060 221.600 151.560 221.700 ;
        RECT 98.550 221.300 151.560 221.600 ;
        RECT 50.680 221.250 51.080 221.300 ;
        RECT 98.550 221.275 98.950 221.300 ;
        RECT 81.150 221.000 81.650 221.100 ;
        RECT 154.740 221.000 155.240 221.100 ;
        RECT 62.640 220.700 81.650 221.000 ;
        RECT 110.500 220.700 155.240 221.000 ;
        RECT 62.640 220.650 63.040 220.700 ;
        RECT 110.500 220.625 110.900 220.700 ;
        RECT 84.800 220.400 85.300 220.500 ;
        RECT 74.600 220.100 85.300 220.400 ;
        RECT 74.600 220.050 75.000 220.100 ;
        RECT 86.560 219.800 86.960 219.825 ;
        RECT 88.500 219.800 89.000 219.900 ;
        RECT 11.140 219.645 13.140 219.795 ;
        RECT 14.385 219.645 14.715 219.660 ;
        RECT 11.140 219.345 14.715 219.645 ;
        RECT 86.560 219.500 89.000 219.800 ;
        RECT 144.105 219.645 144.435 219.660 ;
        RECT 148.440 219.645 150.440 219.795 ;
        RECT 86.560 219.475 86.960 219.500 ;
        RECT 11.140 219.195 13.140 219.345 ;
        RECT 14.385 219.330 14.715 219.345 ;
        RECT 144.105 219.345 150.440 219.645 ;
        RECT 144.105 219.330 144.435 219.345 ;
        RECT 148.440 219.195 150.440 219.345 ;
        RECT 11.140 218.285 13.140 218.435 ;
        RECT 13.925 218.285 14.255 218.300 ;
        RECT 11.140 217.985 14.255 218.285 ;
        RECT 11.140 217.835 13.140 217.985 ;
        RECT 13.925 217.970 14.255 217.985 ;
        RECT 145.485 218.285 145.815 218.300 ;
        RECT 148.440 218.285 150.440 218.435 ;
        RECT 145.485 217.985 150.440 218.285 ;
        RECT 145.485 217.970 145.815 217.985 ;
        RECT 32.690 217.630 34.270 217.960 ;
        RECT 148.440 217.835 150.440 217.985 ;
        RECT 40.605 217.605 40.935 217.620 ;
        RECT 139.505 217.605 139.835 217.620 ;
        RECT 40.605 217.305 139.835 217.605 ;
        RECT 40.605 217.290 40.935 217.305 ;
        RECT 139.505 217.290 139.835 217.305 ;
        RECT 11.140 216.925 13.140 217.075 ;
        RECT 17.605 216.925 17.935 216.940 ;
        RECT 11.140 216.625 17.935 216.925 ;
        RECT 11.140 216.475 13.140 216.625 ;
        RECT 17.605 216.610 17.935 216.625 ;
        RECT 21.285 216.925 21.615 216.940 ;
        RECT 91.205 216.925 91.535 216.940 ;
        RECT 21.285 216.625 91.535 216.925 ;
        RECT 21.285 216.610 21.615 216.625 ;
        RECT 91.205 216.610 91.535 216.625 ;
        RECT 141.805 216.925 142.135 216.940 ;
        RECT 148.440 216.925 150.440 217.075 ;
        RECT 141.805 216.625 150.440 216.925 ;
        RECT 141.805 216.610 142.135 216.625 ;
        RECT 148.440 216.475 150.440 216.625 ;
        RECT 24.965 216.245 25.295 216.260 ;
        RECT 46.125 216.245 46.455 216.260 ;
        RECT 55.325 216.245 55.655 216.260 ;
        RECT 24.965 215.945 55.655 216.245 ;
        RECT 24.965 215.930 25.295 215.945 ;
        RECT 46.125 215.930 46.455 215.945 ;
        RECT 55.325 215.930 55.655 215.945 ;
        RECT 65.445 216.245 65.775 216.260 ;
        RECT 135.365 216.245 135.695 216.260 ;
        RECT 65.445 215.945 135.695 216.245 ;
        RECT 65.445 215.930 65.775 215.945 ;
        RECT 135.365 215.930 135.695 215.945 ;
        RECT 11.140 215.565 13.140 215.715 ;
        RECT 15.765 215.565 16.095 215.580 ;
        RECT 11.140 215.265 16.095 215.565 ;
        RECT 11.140 215.115 13.140 215.265 ;
        RECT 15.765 215.250 16.095 215.265 ;
        RECT 37.845 215.565 38.175 215.580 ;
        RECT 117.425 215.565 117.755 215.580 ;
        RECT 37.845 215.265 117.755 215.565 ;
        RECT 37.845 215.250 38.175 215.265 ;
        RECT 117.425 215.250 117.755 215.265 ;
        RECT 145.945 215.565 146.275 215.580 ;
        RECT 148.440 215.565 150.440 215.715 ;
        RECT 145.945 215.265 150.440 215.565 ;
        RECT 145.945 215.250 146.275 215.265 ;
        RECT 29.390 214.910 30.970 215.240 ;
        RECT 148.440 215.115 150.440 215.265 ;
        RECT 68.665 214.885 68.995 214.900 ;
        RECT 79.245 214.885 79.575 214.900 ;
        RECT 85.685 214.885 86.015 214.900 ;
        RECT 68.665 214.585 86.015 214.885 ;
        RECT 68.665 214.570 68.995 214.585 ;
        RECT 79.245 214.570 79.575 214.585 ;
        RECT 85.685 214.570 86.015 214.585 ;
        RECT 91.665 214.885 91.995 214.900 ;
        RECT 144.565 214.885 144.895 214.900 ;
        RECT 91.665 214.585 144.895 214.885 ;
        RECT 91.665 214.570 91.995 214.585 ;
        RECT 144.565 214.570 144.895 214.585 ;
        RECT 11.140 214.205 13.140 214.355 ;
        RECT 20.365 214.205 20.695 214.220 ;
        RECT 11.140 213.905 20.695 214.205 ;
        RECT 11.140 213.755 13.140 213.905 ;
        RECT 20.365 213.890 20.695 213.905 ;
        RECT 21.745 214.205 22.075 214.220 ;
        RECT 90.285 214.205 90.615 214.220 ;
        RECT 21.745 213.905 90.615 214.205 ;
        RECT 21.745 213.890 22.075 213.905 ;
        RECT 90.285 213.890 90.615 213.905 ;
        RECT 97.645 214.205 97.975 214.220 ;
        RECT 120.185 214.205 120.515 214.220 ;
        RECT 97.645 213.905 120.515 214.205 ;
        RECT 97.645 213.890 97.975 213.905 ;
        RECT 120.185 213.890 120.515 213.905 ;
        RECT 143.645 214.205 143.975 214.220 ;
        RECT 148.440 214.205 150.440 214.355 ;
        RECT 143.645 213.905 150.440 214.205 ;
        RECT 143.645 213.890 143.975 213.905 ;
        RECT 148.440 213.755 150.440 213.905 ;
        RECT 20.365 213.525 20.695 213.540 ;
        RECT 71.425 213.525 71.755 213.540 ;
        RECT 20.365 213.225 71.755 213.525 ;
        RECT 20.365 213.210 20.695 213.225 ;
        RECT 71.425 213.210 71.755 213.225 ;
        RECT 72.345 213.525 72.675 213.540 ;
        RECT 86.145 213.525 86.475 213.540 ;
        RECT 72.345 213.225 86.475 213.525 ;
        RECT 72.345 213.210 72.675 213.225 ;
        RECT 86.145 213.210 86.475 213.225 ;
        RECT 87.065 213.525 87.395 213.540 ;
        RECT 101.785 213.525 102.115 213.540 ;
        RECT 87.065 213.225 102.115 213.525 ;
        RECT 87.065 213.210 87.395 213.225 ;
        RECT 101.785 213.210 102.115 213.225 ;
        RECT 11.140 212.845 13.140 212.995 ;
        RECT 14.845 212.845 15.175 212.860 ;
        RECT 11.140 212.545 15.175 212.845 ;
        RECT 11.140 212.395 13.140 212.545 ;
        RECT 14.845 212.530 15.175 212.545 ;
        RECT 62.225 212.845 62.555 212.860 ;
        RECT 102.245 212.845 102.575 212.860 ;
        RECT 113.285 212.845 113.615 212.860 ;
        RECT 62.225 212.545 113.615 212.845 ;
        RECT 62.225 212.530 62.555 212.545 ;
        RECT 102.245 212.530 102.575 212.545 ;
        RECT 113.285 212.530 113.615 212.545 ;
        RECT 145.485 212.845 145.815 212.860 ;
        RECT 148.440 212.845 150.440 212.995 ;
        RECT 145.485 212.545 150.440 212.845 ;
        RECT 145.485 212.530 145.815 212.545 ;
        RECT 32.690 212.190 34.270 212.520 ;
        RECT 148.440 212.395 150.440 212.545 ;
        RECT 41.065 212.165 41.395 212.180 ;
        RECT 77.865 212.165 78.195 212.180 ;
        RECT 41.065 211.865 78.195 212.165 ;
        RECT 41.065 211.850 41.395 211.865 ;
        RECT 77.865 211.850 78.195 211.865 ;
        RECT 97.185 212.165 97.515 212.180 ;
        RECT 108.225 212.165 108.555 212.180 ;
        RECT 136.745 212.165 137.075 212.180 ;
        RECT 140.885 212.165 141.215 212.180 ;
        RECT 97.185 211.865 141.215 212.165 ;
        RECT 97.185 211.850 97.515 211.865 ;
        RECT 108.225 211.850 108.555 211.865 ;
        RECT 136.745 211.850 137.075 211.865 ;
        RECT 140.885 211.850 141.215 211.865 ;
        RECT 11.140 211.485 13.140 211.635 ;
        RECT 14.385 211.485 14.715 211.500 ;
        RECT 11.140 211.185 14.715 211.485 ;
        RECT 11.140 211.035 13.140 211.185 ;
        RECT 14.385 211.170 14.715 211.185 ;
        RECT 25.425 211.485 25.755 211.500 ;
        RECT 26.805 211.485 27.135 211.500 ;
        RECT 37.385 211.485 37.715 211.500 ;
        RECT 25.425 211.185 37.715 211.485 ;
        RECT 25.425 211.170 25.755 211.185 ;
        RECT 26.805 211.170 27.135 211.185 ;
        RECT 37.385 211.170 37.715 211.185 ;
        RECT 54.865 211.485 55.195 211.500 ;
        RECT 79.705 211.485 80.035 211.500 ;
        RECT 82.005 211.485 82.335 211.500 ;
        RECT 139.045 211.485 139.375 211.500 ;
        RECT 54.865 211.185 139.375 211.485 ;
        RECT 54.865 211.170 55.195 211.185 ;
        RECT 79.705 211.170 80.035 211.185 ;
        RECT 82.005 211.170 82.335 211.185 ;
        RECT 139.045 211.170 139.375 211.185 ;
        RECT 145.485 211.485 145.815 211.500 ;
        RECT 148.440 211.485 150.440 211.635 ;
        RECT 145.485 211.185 150.440 211.485 ;
        RECT 145.485 211.170 145.815 211.185 ;
        RECT 148.440 211.035 150.440 211.185 ;
        RECT 36.925 210.805 37.255 210.820 ;
        RECT 78.785 210.805 79.115 210.820 ;
        RECT 112.825 210.805 113.155 210.820 ;
        RECT 36.925 210.505 113.155 210.805 ;
        RECT 36.925 210.490 37.255 210.505 ;
        RECT 78.785 210.490 79.115 210.505 ;
        RECT 112.825 210.490 113.155 210.505 ;
        RECT 11.140 210.125 13.140 210.275 ;
        RECT 14.505 210.125 14.835 210.140 ;
        RECT 11.140 209.825 14.835 210.125 ;
        RECT 11.140 209.675 13.140 209.825 ;
        RECT 14.505 209.810 14.835 209.825 ;
        RECT 41.525 210.125 41.855 210.140 ;
        RECT 56.245 210.125 56.575 210.140 ;
        RECT 41.525 209.825 56.575 210.125 ;
        RECT 41.525 209.810 41.855 209.825 ;
        RECT 56.245 209.810 56.575 209.825 ;
        RECT 72.345 210.125 72.675 210.140 ;
        RECT 74.645 210.125 74.975 210.140 ;
        RECT 72.345 209.825 74.975 210.125 ;
        RECT 72.345 209.810 72.675 209.825 ;
        RECT 74.645 209.810 74.975 209.825 ;
        RECT 114.205 210.125 114.535 210.140 ;
        RECT 127.545 210.125 127.875 210.140 ;
        RECT 114.205 209.825 127.875 210.125 ;
        RECT 114.205 209.810 114.535 209.825 ;
        RECT 127.545 209.810 127.875 209.825 ;
        RECT 141.805 210.125 142.135 210.140 ;
        RECT 148.440 210.125 150.440 210.275 ;
        RECT 141.805 209.825 150.440 210.125 ;
        RECT 141.805 209.810 142.135 209.825 ;
        RECT 29.390 209.470 30.970 209.800 ;
        RECT 148.440 209.675 150.440 209.825 ;
        RECT 54.865 209.445 55.195 209.460 ;
        RECT 49.130 209.145 55.195 209.445 ;
        RECT 11.140 208.765 13.140 208.915 ;
        RECT 14.165 208.765 14.495 208.780 ;
        RECT 11.140 208.465 14.495 208.765 ;
        RECT 11.140 208.315 13.140 208.465 ;
        RECT 14.165 208.450 14.495 208.465 ;
        RECT 18.525 208.765 18.855 208.780 ;
        RECT 49.130 208.765 49.430 209.145 ;
        RECT 54.865 209.130 55.195 209.145 ;
        RECT 70.505 209.445 70.835 209.460 ;
        RECT 76.025 209.445 76.355 209.460 ;
        RECT 144.565 209.445 144.895 209.460 ;
        RECT 70.505 209.145 144.895 209.445 ;
        RECT 70.505 209.130 70.835 209.145 ;
        RECT 76.025 209.130 76.355 209.145 ;
        RECT 144.565 209.130 144.895 209.145 ;
        RECT 18.525 208.465 49.430 208.765 ;
        RECT 50.265 208.765 50.595 208.780 ;
        RECT 96.265 208.765 96.595 208.780 ;
        RECT 105.005 208.765 105.335 208.780 ;
        RECT 50.265 208.465 91.290 208.765 ;
        RECT 18.525 208.450 18.855 208.465 ;
        RECT 50.265 208.450 50.595 208.465 ;
        RECT 16.685 208.085 17.015 208.100 ;
        RECT 53.025 208.085 53.355 208.100 ;
        RECT 16.685 207.785 53.355 208.085 ;
        RECT 90.990 208.085 91.290 208.465 ;
        RECT 96.265 208.465 105.335 208.765 ;
        RECT 96.265 208.450 96.595 208.465 ;
        RECT 105.005 208.450 105.335 208.465 ;
        RECT 106.385 208.765 106.715 208.780 ;
        RECT 118.805 208.765 119.135 208.780 ;
        RECT 106.385 208.465 119.135 208.765 ;
        RECT 106.385 208.450 106.715 208.465 ;
        RECT 118.805 208.450 119.135 208.465 ;
        RECT 143.645 208.765 143.975 208.780 ;
        RECT 148.440 208.765 150.440 208.915 ;
        RECT 143.645 208.465 150.440 208.765 ;
        RECT 143.645 208.450 143.975 208.465 ;
        RECT 148.440 208.315 150.440 208.465 ;
        RECT 100.865 208.085 101.195 208.100 ;
        RECT 110.065 208.085 110.395 208.100 ;
        RECT 90.990 207.785 110.395 208.085 ;
        RECT 16.685 207.770 17.015 207.785 ;
        RECT 53.025 207.770 53.355 207.785 ;
        RECT 100.865 207.770 101.195 207.785 ;
        RECT 110.065 207.770 110.395 207.785 ;
        RECT 112.365 208.085 112.695 208.100 ;
        RECT 115.585 208.085 115.915 208.100 ;
        RECT 128.925 208.085 129.255 208.100 ;
        RECT 112.365 207.785 129.255 208.085 ;
        RECT 112.365 207.770 112.695 207.785 ;
        RECT 115.585 207.770 115.915 207.785 ;
        RECT 128.925 207.770 129.255 207.785 ;
        RECT 11.140 207.405 13.140 207.555 ;
        RECT 17.605 207.405 17.935 207.420 ;
        RECT 11.140 207.105 17.935 207.405 ;
        RECT 11.140 206.955 13.140 207.105 ;
        RECT 17.605 207.090 17.935 207.105 ;
        RECT 45.205 207.405 45.535 207.420 ;
        RECT 50.265 207.405 50.595 207.420 ;
        RECT 45.205 207.105 50.595 207.405 ;
        RECT 45.205 207.090 45.535 207.105 ;
        RECT 50.265 207.090 50.595 207.105 ;
        RECT 82.925 207.405 83.255 207.420 ;
        RECT 87.065 207.405 87.395 207.420 ;
        RECT 82.925 207.105 87.395 207.405 ;
        RECT 82.925 207.090 83.255 207.105 ;
        RECT 87.065 207.090 87.395 207.105 ;
        RECT 93.505 207.405 93.835 207.420 ;
        RECT 97.645 207.405 97.975 207.420 ;
        RECT 105.465 207.415 105.795 207.420 ;
        RECT 105.210 207.405 105.795 207.415 ;
        RECT 93.505 207.105 97.975 207.405 ;
        RECT 105.010 207.105 105.795 207.405 ;
        RECT 93.505 207.090 93.835 207.105 ;
        RECT 97.645 207.090 97.975 207.105 ;
        RECT 105.210 207.095 105.795 207.105 ;
        RECT 105.465 207.090 105.795 207.095 ;
        RECT 145.485 207.405 145.815 207.420 ;
        RECT 148.440 207.405 150.440 207.555 ;
        RECT 145.485 207.105 150.440 207.405 ;
        RECT 145.485 207.090 145.815 207.105 ;
        RECT 32.690 206.750 34.270 207.080 ;
        RECT 148.440 206.955 150.440 207.105 ;
        RECT 30.485 206.725 30.815 206.740 ;
        RECT 31.610 206.725 31.990 206.735 ;
        RECT 30.485 206.425 31.990 206.725 ;
        RECT 30.485 206.410 30.815 206.425 ;
        RECT 31.610 206.415 31.990 206.425 ;
        RECT 76.485 206.725 76.815 206.740 ;
        RECT 102.705 206.725 103.035 206.740 ;
        RECT 76.485 206.425 103.035 206.725 ;
        RECT 76.485 206.410 76.815 206.425 ;
        RECT 102.705 206.410 103.035 206.425 ;
        RECT 103.625 206.725 103.955 206.740 ;
        RECT 142.725 206.725 143.055 206.740 ;
        RECT 103.625 206.425 143.055 206.725 ;
        RECT 103.625 206.410 103.955 206.425 ;
        RECT 142.725 206.410 143.055 206.425 ;
        RECT 11.140 206.045 13.140 206.195 ;
        RECT 14.085 206.045 14.415 206.060 ;
        RECT 11.140 205.745 14.415 206.045 ;
        RECT 11.140 205.595 13.140 205.745 ;
        RECT 14.085 205.730 14.415 205.745 ;
        RECT 19.445 206.045 19.775 206.060 ;
        RECT 46.125 206.045 46.455 206.060 ;
        RECT 19.445 205.745 46.455 206.045 ;
        RECT 19.445 205.730 19.775 205.745 ;
        RECT 46.125 205.730 46.455 205.745 ;
        RECT 47.045 206.045 47.375 206.060 ;
        RECT 49.805 206.045 50.135 206.060 ;
        RECT 47.045 205.745 50.135 206.045 ;
        RECT 47.045 205.730 47.375 205.745 ;
        RECT 49.805 205.730 50.135 205.745 ;
        RECT 53.945 206.045 54.275 206.060 ;
        RECT 55.785 206.045 56.115 206.060 ;
        RECT 57.165 206.045 57.495 206.060 ;
        RECT 53.945 205.745 57.495 206.045 ;
        RECT 53.945 205.730 54.275 205.745 ;
        RECT 55.785 205.730 56.115 205.745 ;
        RECT 57.165 205.730 57.495 205.745 ;
        RECT 62.225 206.045 62.555 206.060 ;
        RECT 89.365 206.045 89.695 206.060 ;
        RECT 113.285 206.045 113.615 206.060 ;
        RECT 62.225 205.745 113.615 206.045 ;
        RECT 62.225 205.730 62.555 205.745 ;
        RECT 89.365 205.730 89.695 205.745 ;
        RECT 113.285 205.730 113.615 205.745 ;
        RECT 141.805 206.045 142.135 206.060 ;
        RECT 148.440 206.045 150.440 206.195 ;
        RECT 141.805 205.745 150.440 206.045 ;
        RECT 141.805 205.730 142.135 205.745 ;
        RECT 148.440 205.595 150.440 205.745 ;
        RECT 17.145 205.365 17.475 205.380 ;
        RECT 86.605 205.365 86.935 205.380 ;
        RECT 17.145 205.065 86.935 205.365 ;
        RECT 17.145 205.050 17.475 205.065 ;
        RECT 86.605 205.050 86.935 205.065 ;
        RECT 113.745 205.365 114.075 205.380 ;
        RECT 131.685 205.365 132.015 205.380 ;
        RECT 113.745 205.065 132.015 205.365 ;
        RECT 113.745 205.050 114.075 205.065 ;
        RECT 131.685 205.050 132.015 205.065 ;
        RECT 11.140 204.685 13.140 204.835 ;
        RECT 14.055 204.685 14.385 204.700 ;
        RECT 11.140 204.385 14.385 204.685 ;
        RECT 11.140 204.235 13.140 204.385 ;
        RECT 14.055 204.370 14.385 204.385 ;
        RECT 32.785 204.685 33.115 204.700 ;
        RECT 45.665 204.685 45.995 204.700 ;
        RECT 32.785 204.385 45.995 204.685 ;
        RECT 32.785 204.370 33.115 204.385 ;
        RECT 45.665 204.370 45.995 204.385 ;
        RECT 87.065 204.685 87.395 204.700 ;
        RECT 121.105 204.685 121.435 204.700 ;
        RECT 87.065 204.385 121.435 204.685 ;
        RECT 87.065 204.370 87.395 204.385 ;
        RECT 121.105 204.370 121.435 204.385 ;
        RECT 145.485 204.685 145.815 204.700 ;
        RECT 148.440 204.685 150.440 204.835 ;
        RECT 145.485 204.385 150.440 204.685 ;
        RECT 145.485 204.370 145.815 204.385 ;
        RECT 29.390 204.030 30.970 204.360 ;
        RECT 148.440 204.235 150.440 204.385 ;
        RECT 58.085 204.005 58.415 204.020 ;
        RECT 72.345 204.005 72.675 204.020 ;
        RECT 58.085 203.705 72.675 204.005 ;
        RECT 58.085 203.690 58.415 203.705 ;
        RECT 72.345 203.690 72.675 203.705 ;
        RECT 73.725 204.005 74.055 204.020 ;
        RECT 114.205 204.005 114.535 204.020 ;
        RECT 73.725 203.705 114.535 204.005 ;
        RECT 73.725 203.690 74.055 203.705 ;
        RECT 114.205 203.690 114.535 203.705 ;
        RECT 11.140 203.325 13.140 203.475 ;
        RECT 13.925 203.325 14.255 203.340 ;
        RECT 11.140 203.025 14.255 203.325 ;
        RECT 11.140 202.875 13.140 203.025 ;
        RECT 13.925 203.010 14.255 203.025 ;
        RECT 16.685 203.325 17.015 203.340 ;
        RECT 87.525 203.325 87.855 203.340 ;
        RECT 16.685 203.025 87.855 203.325 ;
        RECT 16.685 203.010 17.015 203.025 ;
        RECT 87.525 203.010 87.855 203.025 ;
        RECT 93.505 203.325 93.835 203.340 ;
        RECT 113.745 203.325 114.075 203.340 ;
        RECT 93.505 203.025 114.075 203.325 ;
        RECT 93.505 203.010 93.835 203.025 ;
        RECT 113.745 203.010 114.075 203.025 ;
        RECT 122.945 203.325 123.275 203.340 ;
        RECT 125.245 203.325 125.575 203.340 ;
        RECT 129.845 203.325 130.175 203.340 ;
        RECT 122.945 203.025 130.175 203.325 ;
        RECT 122.945 203.010 123.275 203.025 ;
        RECT 125.245 203.010 125.575 203.025 ;
        RECT 129.845 203.010 130.175 203.025 ;
        RECT 141.805 203.325 142.135 203.340 ;
        RECT 148.440 203.325 150.440 203.475 ;
        RECT 141.805 203.025 150.440 203.325 ;
        RECT 141.805 203.010 142.135 203.025 ;
        RECT 148.440 202.875 150.440 203.025 ;
        RECT 18.065 202.645 18.395 202.660 ;
        RECT 92.125 202.645 92.455 202.660 ;
        RECT 18.065 202.345 92.455 202.645 ;
        RECT 18.065 202.330 18.395 202.345 ;
        RECT 92.125 202.330 92.455 202.345 ;
        RECT 93.965 202.645 94.295 202.660 ;
        RECT 101.325 202.645 101.655 202.660 ;
        RECT 93.965 202.345 101.655 202.645 ;
        RECT 93.965 202.330 94.295 202.345 ;
        RECT 101.325 202.330 101.655 202.345 ;
        RECT 103.165 202.645 103.495 202.660 ;
        RECT 104.085 202.645 104.415 202.660 ;
        RECT 103.165 202.345 104.415 202.645 ;
        RECT 103.165 202.330 103.495 202.345 ;
        RECT 104.085 202.330 104.415 202.345 ;
        RECT 106.845 202.645 107.175 202.660 ;
        RECT 114.665 202.645 114.995 202.660 ;
        RECT 106.845 202.345 114.995 202.645 ;
        RECT 106.845 202.330 107.175 202.345 ;
        RECT 114.665 202.330 114.995 202.345 ;
        RECT 11.140 201.965 13.140 202.115 ;
        RECT 15.765 201.965 16.095 201.980 ;
        RECT 11.140 201.665 16.095 201.965 ;
        RECT 11.140 201.515 13.140 201.665 ;
        RECT 15.765 201.650 16.095 201.665 ;
        RECT 47.965 201.965 48.295 201.980 ;
        RECT 51.850 201.965 52.230 201.975 ;
        RECT 47.965 201.665 52.230 201.965 ;
        RECT 47.965 201.650 48.295 201.665 ;
        RECT 51.850 201.655 52.230 201.665 ;
        RECT 89.365 201.965 89.695 201.980 ;
        RECT 140.885 201.965 141.215 201.980 ;
        RECT 89.365 201.665 141.215 201.965 ;
        RECT 89.365 201.650 89.695 201.665 ;
        RECT 140.885 201.650 141.215 201.665 ;
        RECT 143.645 201.965 143.975 201.980 ;
        RECT 148.440 201.965 150.440 202.115 ;
        RECT 143.645 201.665 150.440 201.965 ;
        RECT 143.645 201.650 143.975 201.665 ;
        RECT 32.690 201.310 34.270 201.640 ;
        RECT 148.440 201.515 150.440 201.665 ;
        RECT 35.545 201.285 35.875 201.300 ;
        RECT 35.330 200.970 35.875 201.285 ;
        RECT 50.265 201.285 50.595 201.300 ;
        RECT 56.705 201.285 57.035 201.300 ;
        RECT 76.945 201.285 77.275 201.300 ;
        RECT 97.185 201.285 97.515 201.300 ;
        RECT 50.265 200.985 97.515 201.285 ;
        RECT 50.265 200.970 50.595 200.985 ;
        RECT 56.705 200.970 57.035 200.985 ;
        RECT 76.945 200.970 77.275 200.985 ;
        RECT 97.185 200.970 97.515 200.985 ;
        RECT 98.105 201.285 98.435 201.300 ;
        RECT 102.705 201.285 103.035 201.300 ;
        RECT 98.105 200.985 103.035 201.285 ;
        RECT 98.105 200.970 98.435 200.985 ;
        RECT 102.705 200.970 103.035 200.985 ;
        RECT 109.605 201.285 109.935 201.300 ;
        RECT 114.205 201.285 114.535 201.300 ;
        RECT 109.605 200.985 114.535 201.285 ;
        RECT 109.605 200.970 109.935 200.985 ;
        RECT 114.205 200.970 114.535 200.985 ;
        RECT 11.140 200.605 13.140 200.755 ;
        RECT 17.605 200.605 17.935 200.620 ;
        RECT 11.140 200.305 17.935 200.605 ;
        RECT 11.140 200.155 13.140 200.305 ;
        RECT 17.605 200.290 17.935 200.305 ;
        RECT 33.705 200.605 34.035 200.620 ;
        RECT 35.330 200.605 35.630 200.970 ;
        RECT 90.745 200.605 91.075 200.620 ;
        RECT 33.705 200.305 35.630 200.605 ;
        RECT 42.690 200.305 91.075 200.605 ;
        RECT 33.705 200.290 34.035 200.305 ;
        RECT 16.685 199.925 17.015 199.940 ;
        RECT 42.690 199.925 42.990 200.305 ;
        RECT 90.745 200.290 91.075 200.305 ;
        RECT 93.045 200.605 93.375 200.620 ;
        RECT 109.605 200.605 109.935 200.620 ;
        RECT 128.465 200.605 128.795 200.620 ;
        RECT 131.685 200.605 132.015 200.620 ;
        RECT 132.605 200.605 132.935 200.620 ;
        RECT 93.045 200.305 132.935 200.605 ;
        RECT 93.045 200.290 93.375 200.305 ;
        RECT 109.605 200.290 109.935 200.305 ;
        RECT 128.465 200.290 128.795 200.305 ;
        RECT 131.685 200.290 132.015 200.305 ;
        RECT 132.605 200.290 132.935 200.305 ;
        RECT 145.485 200.605 145.815 200.620 ;
        RECT 148.440 200.605 150.440 200.755 ;
        RECT 145.485 200.305 150.440 200.605 ;
        RECT 145.485 200.290 145.815 200.305 ;
        RECT 148.440 200.155 150.440 200.305 ;
        RECT 16.685 199.625 42.990 199.925 ;
        RECT 45.205 199.925 45.535 199.940 ;
        RECT 52.565 199.925 52.895 199.940 ;
        RECT 45.205 199.625 52.895 199.925 ;
        RECT 16.685 199.610 17.015 199.625 ;
        RECT 45.205 199.610 45.535 199.625 ;
        RECT 52.565 199.610 52.895 199.625 ;
        RECT 56.705 199.925 57.035 199.940 ;
        RECT 59.925 199.925 60.255 199.940 ;
        RECT 110.985 199.925 111.315 199.940 ;
        RECT 56.705 199.625 111.315 199.925 ;
        RECT 56.705 199.610 57.035 199.625 ;
        RECT 59.925 199.610 60.255 199.625 ;
        RECT 110.985 199.610 111.315 199.625 ;
        RECT 112.825 199.925 113.155 199.940 ;
        RECT 128.465 199.925 128.795 199.940 ;
        RECT 112.825 199.625 128.795 199.925 ;
        RECT 112.825 199.610 113.155 199.625 ;
        RECT 128.465 199.610 128.795 199.625 ;
        RECT 11.140 199.245 13.140 199.395 ;
        RECT 14.845 199.245 15.175 199.260 ;
        RECT 11.140 198.945 15.175 199.245 ;
        RECT 11.140 198.795 13.140 198.945 ;
        RECT 14.845 198.930 15.175 198.945 ;
        RECT 34.165 199.245 34.495 199.260 ;
        RECT 40.145 199.245 40.475 199.260 ;
        RECT 44.285 199.245 44.615 199.260 ;
        RECT 50.265 199.245 50.595 199.260 ;
        RECT 34.165 198.945 50.595 199.245 ;
        RECT 34.165 198.930 34.495 198.945 ;
        RECT 40.145 198.930 40.475 198.945 ;
        RECT 44.285 198.930 44.615 198.945 ;
        RECT 50.265 198.930 50.595 198.945 ;
        RECT 54.405 199.245 54.735 199.260 ;
        RECT 67.285 199.245 67.615 199.260 ;
        RECT 82.925 199.245 83.255 199.260 ;
        RECT 54.405 198.945 83.255 199.245 ;
        RECT 54.405 198.930 54.735 198.945 ;
        RECT 67.285 198.930 67.615 198.945 ;
        RECT 82.925 198.930 83.255 198.945 ;
        RECT 87.065 199.245 87.395 199.260 ;
        RECT 140.885 199.245 141.215 199.260 ;
        RECT 87.065 198.945 141.215 199.245 ;
        RECT 87.065 198.930 87.395 198.945 ;
        RECT 140.885 198.930 141.215 198.945 ;
        RECT 145.485 199.245 145.815 199.260 ;
        RECT 148.440 199.245 150.440 199.395 ;
        RECT 145.485 198.945 150.440 199.245 ;
        RECT 145.485 198.930 145.815 198.945 ;
        RECT 29.390 198.590 30.970 198.920 ;
        RECT 148.440 198.795 150.440 198.945 ;
        RECT 24.505 198.565 24.835 198.580 ;
        RECT 26.345 198.565 26.675 198.580 ;
        RECT 24.505 198.265 26.675 198.565 ;
        RECT 24.505 198.250 24.835 198.265 ;
        RECT 26.345 198.250 26.675 198.265 ;
        RECT 32.325 198.565 32.655 198.580 ;
        RECT 44.745 198.565 45.075 198.580 ;
        RECT 32.325 198.265 45.075 198.565 ;
        RECT 32.325 198.250 32.655 198.265 ;
        RECT 44.745 198.250 45.075 198.265 ;
        RECT 50.265 198.565 50.595 198.580 ;
        RECT 57.625 198.565 57.955 198.580 ;
        RECT 59.465 198.565 59.795 198.580 ;
        RECT 50.265 198.265 59.795 198.565 ;
        RECT 50.265 198.250 50.595 198.265 ;
        RECT 57.625 198.250 57.955 198.265 ;
        RECT 59.465 198.250 59.795 198.265 ;
        RECT 95.345 198.565 95.675 198.580 ;
        RECT 100.405 198.565 100.735 198.580 ;
        RECT 95.345 198.265 100.735 198.565 ;
        RECT 95.345 198.250 95.675 198.265 ;
        RECT 100.405 198.250 100.735 198.265 ;
        RECT 101.325 198.565 101.655 198.580 ;
        RECT 132.605 198.565 132.935 198.580 ;
        RECT 101.325 198.265 132.935 198.565 ;
        RECT 101.325 198.250 101.655 198.265 ;
        RECT 132.605 198.250 132.935 198.265 ;
        RECT 11.140 197.885 13.140 198.035 ;
        RECT 14.385 197.885 14.715 197.900 ;
        RECT 11.140 197.585 14.715 197.885 ;
        RECT 11.140 197.435 13.140 197.585 ;
        RECT 14.385 197.570 14.715 197.585 ;
        RECT 31.610 197.885 31.990 197.895 ;
        RECT 35.085 197.885 35.415 197.900 ;
        RECT 31.610 197.585 35.415 197.885 ;
        RECT 31.610 197.575 31.990 197.585 ;
        RECT 35.085 197.570 35.415 197.585 ;
        RECT 46.125 197.885 46.455 197.900 ;
        RECT 102.705 197.885 103.035 197.900 ;
        RECT 46.125 197.585 103.035 197.885 ;
        RECT 46.125 197.570 46.455 197.585 ;
        RECT 102.705 197.570 103.035 197.585 ;
        RECT 141.805 197.885 142.135 197.900 ;
        RECT 148.440 197.885 150.440 198.035 ;
        RECT 141.805 197.585 150.440 197.885 ;
        RECT 141.805 197.570 142.135 197.585 ;
        RECT 148.440 197.435 150.440 197.585 ;
        RECT 29.565 197.205 29.895 197.220 ;
        RECT 33.705 197.205 34.035 197.220 ;
        RECT 29.565 196.905 34.035 197.205 ;
        RECT 29.565 196.890 29.895 196.905 ;
        RECT 33.705 196.890 34.035 196.905 ;
        RECT 35.545 197.205 35.875 197.220 ;
        RECT 48.885 197.205 49.215 197.220 ;
        RECT 35.545 196.905 49.215 197.205 ;
        RECT 35.545 196.890 35.875 196.905 ;
        RECT 48.885 196.890 49.215 196.905 ;
        RECT 51.850 197.205 52.230 197.215 ;
        RECT 52.565 197.205 52.895 197.220 ;
        RECT 51.850 196.905 52.895 197.205 ;
        RECT 51.850 196.895 52.230 196.905 ;
        RECT 52.565 196.890 52.895 196.905 ;
        RECT 71.885 197.205 72.215 197.220 ;
        RECT 74.645 197.205 74.975 197.220 ;
        RECT 71.885 196.905 74.975 197.205 ;
        RECT 71.885 196.890 72.215 196.905 ;
        RECT 74.645 196.890 74.975 196.905 ;
        RECT 81.545 197.205 81.875 197.220 ;
        RECT 142.725 197.205 143.055 197.220 ;
        RECT 81.545 196.905 143.055 197.205 ;
        RECT 81.545 196.890 81.875 196.905 ;
        RECT 142.725 196.890 143.055 196.905 ;
        RECT 11.140 196.525 13.140 196.675 ;
        RECT 14.845 196.525 15.175 196.540 ;
        RECT 11.140 196.225 15.175 196.525 ;
        RECT 11.140 196.075 13.140 196.225 ;
        RECT 14.845 196.210 15.175 196.225 ;
        RECT 36.925 196.525 37.255 196.540 ;
        RECT 73.265 196.525 73.595 196.540 ;
        RECT 106.385 196.525 106.715 196.540 ;
        RECT 36.925 196.225 58.630 196.525 ;
        RECT 36.925 196.210 37.255 196.225 ;
        RECT 32.690 195.870 34.270 196.200 ;
        RECT 38.305 195.845 38.635 195.860 ;
        RECT 40.605 195.845 40.935 195.860 ;
        RECT 46.585 195.845 46.915 195.860 ;
        RECT 54.865 195.845 55.195 195.860 ;
        RECT 38.305 195.545 55.195 195.845 ;
        RECT 58.330 195.845 58.630 196.225 ;
        RECT 73.265 196.225 106.715 196.525 ;
        RECT 73.265 196.210 73.595 196.225 ;
        RECT 106.385 196.210 106.715 196.225 ;
        RECT 132.605 196.525 132.935 196.540 ;
        RECT 139.965 196.525 140.295 196.540 ;
        RECT 132.605 196.225 140.295 196.525 ;
        RECT 132.605 196.210 132.935 196.225 ;
        RECT 139.965 196.210 140.295 196.225 ;
        RECT 143.645 196.525 143.975 196.540 ;
        RECT 148.440 196.525 150.440 196.675 ;
        RECT 143.645 196.225 150.440 196.525 ;
        RECT 143.645 196.210 143.975 196.225 ;
        RECT 148.440 196.075 150.440 196.225 ;
        RECT 62.685 195.845 63.015 195.860 ;
        RECT 71.885 195.845 72.215 195.860 ;
        RECT 58.330 195.545 72.215 195.845 ;
        RECT 38.305 195.530 38.635 195.545 ;
        RECT 40.605 195.530 40.935 195.545 ;
        RECT 46.585 195.530 46.915 195.545 ;
        RECT 54.865 195.530 55.195 195.545 ;
        RECT 62.685 195.530 63.015 195.545 ;
        RECT 71.885 195.530 72.215 195.545 ;
        RECT 82.925 195.845 83.255 195.860 ;
        RECT 104.085 195.845 104.415 195.860 ;
        RECT 82.925 195.545 104.415 195.845 ;
        RECT 82.925 195.530 83.255 195.545 ;
        RECT 104.085 195.530 104.415 195.545 ;
        RECT 105.005 195.855 105.335 195.860 ;
        RECT 105.005 195.845 105.590 195.855 ;
        RECT 110.525 195.845 110.855 195.860 ;
        RECT 128.005 195.845 128.335 195.860 ;
        RECT 105.005 195.545 105.790 195.845 ;
        RECT 110.525 195.545 128.335 195.845 ;
        RECT 105.005 195.535 105.590 195.545 ;
        RECT 105.005 195.530 105.335 195.535 ;
        RECT 110.525 195.530 110.855 195.545 ;
        RECT 128.005 195.530 128.335 195.545 ;
        RECT 128.925 195.845 129.255 195.860 ;
        RECT 143.185 195.845 143.515 195.860 ;
        RECT 128.925 195.545 143.515 195.845 ;
        RECT 128.925 195.530 129.255 195.545 ;
        RECT 143.185 195.530 143.515 195.545 ;
        RECT 11.140 195.165 13.140 195.315 ;
        RECT 15.765 195.165 16.095 195.180 ;
        RECT 11.140 194.865 16.095 195.165 ;
        RECT 11.140 194.715 13.140 194.865 ;
        RECT 15.765 194.850 16.095 194.865 ;
        RECT 18.065 195.165 18.395 195.180 ;
        RECT 70.045 195.165 70.375 195.180 ;
        RECT 18.065 194.865 70.375 195.165 ;
        RECT 18.065 194.850 18.395 194.865 ;
        RECT 70.045 194.850 70.375 194.865 ;
        RECT 82.465 195.165 82.795 195.180 ;
        RECT 144.565 195.165 144.895 195.180 ;
        RECT 82.465 194.865 144.895 195.165 ;
        RECT 82.465 194.850 82.795 194.865 ;
        RECT 144.565 194.850 144.895 194.865 ;
        RECT 145.485 195.165 145.815 195.180 ;
        RECT 148.440 195.165 150.440 195.315 ;
        RECT 145.485 194.865 150.440 195.165 ;
        RECT 145.485 194.850 145.815 194.865 ;
        RECT 148.440 194.715 150.440 194.865 ;
        RECT 29.565 194.485 29.895 194.500 ;
        RECT 32.785 194.485 33.115 194.500 ;
        RECT 60.385 194.485 60.715 194.500 ;
        RECT 67.745 194.485 68.075 194.500 ;
        RECT 115.585 194.485 115.915 194.500 ;
        RECT 134.445 194.485 134.775 194.500 ;
        RECT 29.565 194.185 134.775 194.485 ;
        RECT 29.565 194.170 29.895 194.185 ;
        RECT 32.785 194.170 33.115 194.185 ;
        RECT 60.385 194.170 60.715 194.185 ;
        RECT 67.745 194.170 68.075 194.185 ;
        RECT 115.585 194.170 115.915 194.185 ;
        RECT 134.445 194.170 134.775 194.185 ;
        RECT 11.140 193.805 13.140 193.955 ;
        RECT 17.605 193.805 17.935 193.820 ;
        RECT 11.140 193.505 17.935 193.805 ;
        RECT 11.140 193.355 13.140 193.505 ;
        RECT 17.605 193.490 17.935 193.505 ;
        RECT 33.245 193.805 33.575 193.820 ;
        RECT 74.645 193.805 74.975 193.820 ;
        RECT 104.085 193.805 104.415 193.820 ;
        RECT 33.245 193.505 104.415 193.805 ;
        RECT 33.245 193.490 33.575 193.505 ;
        RECT 74.645 193.490 74.975 193.505 ;
        RECT 104.085 193.490 104.415 193.505 ;
        RECT 112.365 193.805 112.695 193.820 ;
        RECT 122.945 193.805 123.275 193.820 ;
        RECT 112.365 193.505 123.275 193.805 ;
        RECT 112.365 193.490 112.695 193.505 ;
        RECT 122.945 193.490 123.275 193.505 ;
        RECT 138.125 193.805 138.455 193.820 ;
        RECT 141.805 193.805 142.135 193.820 ;
        RECT 148.440 193.805 150.440 193.955 ;
        RECT 138.125 193.490 138.670 193.805 ;
        RECT 141.805 193.505 150.440 193.805 ;
        RECT 141.805 193.490 142.135 193.505 ;
        RECT 29.390 193.150 30.970 193.480 ;
        RECT 117.885 193.125 118.215 193.140 ;
        RECT 46.370 192.825 118.215 193.125 ;
        RECT 11.140 192.445 13.140 192.595 ;
        RECT 13.465 192.445 13.795 192.460 ;
        RECT 11.140 192.145 13.795 192.445 ;
        RECT 11.140 191.995 13.140 192.145 ;
        RECT 13.465 192.130 13.795 192.145 ;
        RECT 19.905 192.445 20.235 192.460 ;
        RECT 46.370 192.445 46.670 192.825 ;
        RECT 117.885 192.810 118.215 192.825 ;
        RECT 121.105 193.125 121.435 193.140 ;
        RECT 133.065 193.125 133.395 193.140 ;
        RECT 121.105 192.825 133.395 193.125 ;
        RECT 121.105 192.810 121.435 192.825 ;
        RECT 133.065 192.810 133.395 192.825 ;
        RECT 131.685 192.445 132.015 192.460 ;
        RECT 19.905 192.145 46.670 192.445 ;
        RECT 50.970 192.145 132.015 192.445 ;
        RECT 19.905 192.130 20.235 192.145 ;
        RECT 33.705 191.765 34.035 191.780 ;
        RECT 50.970 191.765 51.270 192.145 ;
        RECT 131.685 192.130 132.015 192.145 ;
        RECT 33.705 191.465 51.270 191.765 ;
        RECT 51.645 191.765 51.975 191.780 ;
        RECT 137.205 191.765 137.535 191.780 ;
        RECT 51.645 191.465 137.535 191.765 ;
        RECT 33.705 191.450 34.035 191.465 ;
        RECT 51.645 191.450 51.975 191.465 ;
        RECT 137.205 191.450 137.535 191.465 ;
        RECT 11.140 191.085 13.140 191.235 ;
        RECT 14.845 191.085 15.175 191.100 ;
        RECT 11.140 190.785 15.175 191.085 ;
        RECT 11.140 190.635 13.140 190.785 ;
        RECT 14.845 190.770 15.175 190.785 ;
        RECT 54.405 191.085 54.735 191.100 ;
        RECT 58.545 191.085 58.875 191.100 ;
        RECT 128.005 191.085 128.335 191.100 ;
        RECT 54.405 190.785 58.875 191.085 ;
        RECT 54.405 190.770 54.735 190.785 ;
        RECT 58.545 190.770 58.875 190.785 ;
        RECT 94.210 190.785 128.335 191.085 ;
        RECT 138.370 191.085 138.670 193.490 ;
        RECT 148.440 193.355 150.440 193.505 ;
        RECT 139.045 192.445 139.375 192.460 ;
        RECT 148.440 192.445 150.440 192.595 ;
        RECT 139.045 192.145 150.440 192.445 ;
        RECT 139.045 192.130 139.375 192.145 ;
        RECT 148.440 191.995 150.440 192.145 ;
        RECT 148.440 191.085 150.440 191.235 ;
        RECT 138.370 190.785 150.440 191.085 ;
        RECT 32.690 190.430 34.270 190.760 ;
        RECT 49.345 190.405 49.675 190.420 ;
        RECT 94.210 190.405 94.510 190.785 ;
        RECT 128.005 190.770 128.335 190.785 ;
        RECT 148.440 190.635 150.440 190.785 ;
        RECT 49.345 190.105 94.510 190.405 ;
        RECT 49.345 190.090 49.675 190.105 ;
        RECT 11.140 189.725 13.140 189.875 ;
        RECT 28.185 189.725 28.515 189.740 ;
        RECT 11.140 189.425 28.515 189.725 ;
        RECT 11.140 189.275 13.140 189.425 ;
        RECT 28.185 189.410 28.515 189.425 ;
        RECT 48.885 189.725 49.215 189.740 ;
        RECT 136.285 189.725 136.615 189.740 ;
        RECT 48.885 189.425 136.615 189.725 ;
        RECT 48.885 189.410 49.215 189.425 ;
        RECT 136.285 189.410 136.615 189.425 ;
        RECT 138.125 189.725 138.455 189.740 ;
        RECT 148.440 189.725 150.440 189.875 ;
        RECT 138.125 189.425 150.440 189.725 ;
        RECT 138.125 189.410 138.455 189.425 ;
        RECT 148.440 189.275 150.440 189.425 ;
        RECT 12.090 189.265 12.490 189.275 ;
        RECT 14.640 183.540 34.390 185.240 ;
        RECT 142.190 184.665 145.090 185.465 ;
        RECT 14.640 182.815 15.490 183.540 ;
        RECT 14.590 182.365 15.540 182.815 ;
        RECT 16.490 182.715 17.340 182.790 ;
        RECT 16.440 182.690 17.390 182.715 ;
        RECT 29.290 182.690 31.090 182.715 ;
        RECT 37.490 182.690 39.440 182.715 ;
        RECT 76.090 182.690 78.040 182.715 ;
        RECT 115.190 182.690 117.140 182.715 ;
        RECT 14.640 177.365 15.490 182.365 ;
        RECT 16.440 180.990 141.790 182.690 ;
        RECT 16.440 180.965 17.390 180.990 ;
        RECT 29.290 180.965 31.090 180.990 ;
        RECT 37.490 180.965 39.440 180.990 ;
        RECT 76.090 180.965 78.040 180.990 ;
        RECT 115.190 180.965 117.140 180.990 ;
        RECT 16.490 180.065 17.340 180.965 ;
        RECT 16.440 179.615 17.390 180.065 ;
        RECT 14.590 176.915 15.540 177.365 ;
        RECT 14.640 171.915 15.490 176.915 ;
        RECT 16.490 174.615 17.340 179.615 ;
        RECT 78.190 178.340 83.290 179.390 ;
        RECT 78.190 176.590 81.040 178.340 ;
        RECT 81.540 177.240 82.040 177.740 ;
        RECT 82.690 176.590 83.290 178.340 ;
        RECT 16.440 174.165 17.390 174.615 ;
        RECT 78.190 174.590 83.290 176.590 ;
        RECT 14.590 171.465 15.540 171.915 ;
        RECT 14.640 166.465 15.490 171.465 ;
        RECT 16.490 169.215 17.340 174.165 ;
        RECT 78.190 172.840 79.040 174.590 ;
        RECT 79.590 173.440 80.140 173.940 ;
        RECT 80.690 172.840 83.290 174.590 ;
        RECT 16.440 168.765 17.390 169.215 ;
        RECT 14.590 166.015 15.540 166.465 ;
        RECT 16.490 166.040 17.340 168.765 ;
        RECT 39.590 165.940 41.390 165.965 ;
        RECT 66.840 165.940 68.640 165.965 ;
        RECT 78.190 165.940 83.290 172.840 ;
        RECT 104.090 168.690 104.490 168.715 ;
        RECT 108.190 168.690 108.590 168.715 ;
        RECT 104.090 168.390 108.590 168.690 ;
        RECT 104.090 168.365 104.490 168.390 ;
        RECT 108.190 168.365 108.590 168.390 ;
        RECT 104.090 168.040 104.490 168.065 ;
        RECT 108.540 168.040 108.940 168.065 ;
        RECT 104.090 167.740 108.940 168.040 ;
        RECT 104.090 167.715 104.490 167.740 ;
        RECT 108.540 167.715 108.940 167.740 ;
        RECT 32.590 164.240 145.090 165.940 ;
        RECT 39.590 164.215 41.390 164.240 ;
        RECT 66.840 164.215 68.640 164.240 ;
        RECT 32.590 159.765 34.390 160.265 ;
        RECT 3.240 157.615 3.640 157.965 ;
        RECT 3.290 135.865 3.590 157.615 ;
        RECT 36.540 157.240 36.940 157.640 ;
        RECT 5.190 153.515 5.590 154.765 ;
        RECT 5.240 140.115 5.540 153.515 ;
        RECT 29.290 152.765 31.090 154.515 ;
        RECT 36.590 153.290 36.890 157.240 ;
        RECT 36.540 152.890 36.940 153.290 ;
        RECT 5.890 141.615 6.190 141.790 ;
        RECT 5.840 141.265 6.240 141.615 ;
        RECT 5.190 139.765 5.590 140.115 ;
        RECT 4.590 138.565 4.890 138.740 ;
        RECT 4.540 138.215 4.940 138.565 ;
        RECT 3.940 136.515 4.240 136.690 ;
        RECT 3.890 136.165 4.290 136.515 ;
        RECT 3.240 135.515 3.640 135.865 ;
        RECT 3.290 2.450 3.590 135.515 ;
        RECT 3.940 3.390 4.240 136.165 ;
        RECT 4.590 4.040 4.890 138.215 ;
        RECT 5.890 137.890 6.190 141.265 ;
        RECT 5.240 137.590 6.190 137.890 ;
        RECT 5.240 4.690 5.540 137.590 ;
        RECT 35.240 133.640 37.040 140.040 ;
        RECT 45.190 139.215 45.590 142.240 ;
        RECT 46.690 141.040 50.790 142.440 ;
        RECT 46.690 139.790 48.190 141.040 ;
        RECT 48.490 140.215 48.990 140.715 ;
        RECT 49.290 139.790 50.790 141.040 ;
        RECT 43.440 136.165 43.840 138.465 ;
        RECT 46.690 133.640 50.790 139.790 ;
        RECT 56.190 135.315 56.590 141.640 ;
        RECT 57.140 138.065 57.540 141.040 ;
        RECT 58.690 134.015 59.090 140.315 ;
        RECT 59.640 134.015 60.040 140.315 ;
        RECT 60.690 134.015 61.090 140.315 ;
        RECT 61.740 134.015 62.140 140.315 ;
        RECT 62.790 134.015 63.190 140.315 ;
        RECT 63.840 134.015 64.240 140.340 ;
        RECT 64.890 134.015 65.290 140.340 ;
        RECT 35.240 133.540 50.790 133.640 ;
        RECT 78.190 133.590 83.290 164.240 ;
        RECT 128.890 160.265 130.590 164.240 ;
        RECT 128.840 159.765 130.640 160.265 ;
        RECT 124.175 157.240 124.575 157.640 ;
        RECT 157.475 157.615 157.875 157.965 ;
        RECT 124.225 153.290 124.525 157.240 ;
        RECT 124.175 152.890 124.575 153.290 ;
        RECT 127.490 152.615 129.440 154.515 ;
        RECT 155.525 153.515 155.925 154.765 ;
        RECT 95.825 134.015 96.225 140.340 ;
        RECT 96.875 134.015 97.275 140.340 ;
        RECT 97.925 134.015 98.325 140.315 ;
        RECT 98.975 134.015 99.375 140.315 ;
        RECT 100.025 134.015 100.425 140.315 ;
        RECT 101.075 134.015 101.475 140.315 ;
        RECT 102.025 134.015 102.425 140.315 ;
        RECT 103.575 138.065 103.975 141.040 ;
        RECT 104.525 135.315 104.925 141.640 ;
        RECT 110.390 141.040 114.490 142.440 ;
        RECT 110.390 139.790 111.790 141.040 ;
        RECT 112.125 140.215 112.625 140.715 ;
        RECT 112.940 139.790 114.490 141.040 ;
        RECT 110.390 133.640 114.490 139.790 ;
        RECT 115.525 139.215 115.925 142.240 ;
        RECT 154.925 141.615 155.225 141.790 ;
        RECT 154.875 141.265 155.275 141.615 ;
        RECT 117.275 136.165 117.675 138.465 ;
        RECT 123.990 138.265 125.890 140.115 ;
        RECT 124.090 133.640 125.890 138.265 ;
        RECT 154.925 137.890 155.225 141.265 ;
        RECT 155.575 140.115 155.875 153.515 ;
        RECT 155.525 139.765 155.925 140.115 ;
        RECT 156.225 138.565 156.525 138.740 ;
        RECT 156.175 138.215 156.575 138.565 ;
        RECT 154.925 137.590 155.875 137.890 ;
        RECT 110.390 133.590 125.890 133.640 ;
        RECT 78.190 133.540 125.890 133.590 ;
        RECT 35.240 131.840 125.890 133.540 ;
        RECT 46.690 129.990 114.490 131.840 ;
        RECT 46.690 129.940 90.890 129.990 ;
        RECT 70.240 128.490 90.890 129.940 ;
        RECT 7.340 127.190 8.340 127.590 ;
        RECT 70.240 126.640 89.890 128.490 ;
        RECT 152.775 127.190 153.775 127.590 ;
        RECT 6.840 125.240 8.540 126.640 ;
        RECT 8.840 125.240 10.540 126.640 ;
        RECT 10.840 125.240 12.540 126.640 ;
        RECT 12.840 125.240 14.540 126.640 ;
        RECT 14.840 125.240 16.540 126.640 ;
        RECT 16.840 125.240 18.540 126.640 ;
        RECT 18.840 125.240 20.540 126.640 ;
        RECT 20.840 125.240 22.540 126.640 ;
        RECT 22.840 125.240 24.540 126.640 ;
        RECT 24.840 125.240 26.540 126.640 ;
        RECT 26.840 125.240 28.540 126.640 ;
        RECT 28.840 125.240 30.540 126.640 ;
        RECT 30.840 125.240 32.540 126.640 ;
        RECT 32.840 125.240 34.540 126.640 ;
        RECT 34.840 125.240 36.540 126.640 ;
        RECT 36.840 125.240 38.540 126.640 ;
        RECT 38.840 125.240 40.540 126.640 ;
        RECT 40.840 125.240 42.540 126.640 ;
        RECT 42.840 125.240 44.540 126.640 ;
        RECT 44.840 125.240 46.540 126.640 ;
        RECT 46.840 125.240 48.540 126.640 ;
        RECT 48.840 125.240 50.540 126.640 ;
        RECT 50.840 125.240 52.540 126.640 ;
        RECT 52.840 125.240 54.540 126.640 ;
        RECT 54.840 125.240 56.540 126.640 ;
        RECT 56.840 125.240 58.540 126.640 ;
        RECT 58.840 125.240 60.540 126.640 ;
        RECT 60.840 125.240 62.540 126.640 ;
        RECT 62.840 125.240 64.540 126.640 ;
        RECT 64.840 125.240 66.540 126.640 ;
        RECT 66.840 125.240 68.540 126.640 ;
        RECT 68.840 125.240 70.540 126.640 ;
        RECT 70.840 125.240 72.540 126.640 ;
        RECT 72.840 125.240 74.540 126.640 ;
        RECT 86.575 125.240 88.275 126.640 ;
        RECT 88.575 125.240 90.275 126.640 ;
        RECT 90.575 125.240 92.275 126.640 ;
        RECT 92.575 125.240 94.275 126.640 ;
        RECT 94.575 125.240 96.275 126.640 ;
        RECT 96.575 125.240 98.275 126.640 ;
        RECT 98.575 125.240 100.275 126.640 ;
        RECT 100.575 125.240 102.275 126.640 ;
        RECT 102.575 125.240 104.275 126.640 ;
        RECT 104.575 125.240 106.275 126.640 ;
        RECT 106.575 125.240 108.275 126.640 ;
        RECT 108.575 125.240 110.275 126.640 ;
        RECT 110.575 125.240 112.275 126.640 ;
        RECT 112.575 125.240 114.275 126.640 ;
        RECT 114.575 125.240 116.275 126.640 ;
        RECT 116.575 125.240 118.275 126.640 ;
        RECT 118.575 125.240 120.275 126.640 ;
        RECT 120.575 125.240 122.275 126.640 ;
        RECT 122.575 125.240 124.275 126.640 ;
        RECT 124.575 125.240 126.275 126.640 ;
        RECT 126.575 125.240 128.275 126.640 ;
        RECT 128.575 125.240 130.275 126.640 ;
        RECT 130.575 125.240 132.275 126.640 ;
        RECT 132.575 125.240 134.275 126.640 ;
        RECT 134.575 125.240 136.275 126.640 ;
        RECT 136.575 125.240 138.275 126.640 ;
        RECT 138.575 125.240 140.275 126.640 ;
        RECT 140.575 125.240 142.275 126.640 ;
        RECT 142.575 125.240 144.275 126.640 ;
        RECT 144.575 125.240 146.275 126.640 ;
        RECT 146.575 125.240 148.275 126.640 ;
        RECT 148.575 125.240 150.275 126.640 ;
        RECT 150.575 125.240 152.275 126.640 ;
        RECT 152.575 125.240 154.275 126.640 ;
        RECT 6.840 123.390 8.540 124.790 ;
        RECT 8.840 123.390 10.540 124.790 ;
        RECT 10.840 123.390 12.540 124.790 ;
        RECT 12.840 123.390 14.540 124.790 ;
        RECT 14.840 123.390 16.540 124.790 ;
        RECT 16.840 123.390 18.540 124.790 ;
        RECT 18.840 123.390 20.540 124.790 ;
        RECT 20.840 123.390 22.540 124.790 ;
        RECT 22.840 123.390 24.540 124.790 ;
        RECT 24.840 123.390 26.540 124.790 ;
        RECT 26.840 123.390 28.540 124.790 ;
        RECT 28.840 123.390 30.540 124.790 ;
        RECT 30.840 123.390 32.540 124.790 ;
        RECT 32.840 123.390 34.540 124.790 ;
        RECT 34.840 123.390 36.540 124.790 ;
        RECT 36.840 123.390 38.540 124.790 ;
        RECT 38.840 123.390 40.540 124.790 ;
        RECT 40.840 123.390 42.540 124.790 ;
        RECT 42.840 123.390 44.540 124.790 ;
        RECT 44.840 123.390 46.540 124.790 ;
        RECT 46.840 123.390 48.540 124.790 ;
        RECT 48.840 123.390 50.540 124.790 ;
        RECT 50.840 123.390 52.540 124.790 ;
        RECT 52.840 123.390 54.540 124.790 ;
        RECT 54.840 123.390 56.540 124.790 ;
        RECT 56.840 123.390 58.540 124.790 ;
        RECT 58.840 123.390 60.540 124.790 ;
        RECT 60.840 123.390 62.540 124.790 ;
        RECT 62.840 123.390 64.540 124.790 ;
        RECT 64.840 123.390 66.540 124.790 ;
        RECT 66.840 123.390 68.540 124.790 ;
        RECT 68.840 123.390 70.540 124.790 ;
        RECT 70.840 123.390 72.540 124.790 ;
        RECT 72.840 123.390 74.540 124.790 ;
        RECT 86.575 123.390 88.275 124.790 ;
        RECT 88.575 123.390 90.275 124.790 ;
        RECT 90.575 123.390 92.275 124.790 ;
        RECT 92.575 123.390 94.275 124.790 ;
        RECT 94.575 123.390 96.275 124.790 ;
        RECT 96.575 123.390 98.275 124.790 ;
        RECT 98.575 123.390 100.275 124.790 ;
        RECT 100.575 123.390 102.275 124.790 ;
        RECT 102.575 123.390 104.275 124.790 ;
        RECT 104.575 123.390 106.275 124.790 ;
        RECT 106.575 123.390 108.275 124.790 ;
        RECT 108.575 123.390 110.275 124.790 ;
        RECT 110.575 123.390 112.275 124.790 ;
        RECT 112.575 123.390 114.275 124.790 ;
        RECT 114.575 123.390 116.275 124.790 ;
        RECT 116.575 123.390 118.275 124.790 ;
        RECT 118.575 123.390 120.275 124.790 ;
        RECT 120.575 123.390 122.275 124.790 ;
        RECT 122.575 123.390 124.275 124.790 ;
        RECT 124.575 123.390 126.275 124.790 ;
        RECT 126.575 123.390 128.275 124.790 ;
        RECT 128.575 123.390 130.275 124.790 ;
        RECT 130.575 123.390 132.275 124.790 ;
        RECT 132.575 123.390 134.275 124.790 ;
        RECT 134.575 123.390 136.275 124.790 ;
        RECT 136.575 123.390 138.275 124.790 ;
        RECT 138.575 123.390 140.275 124.790 ;
        RECT 140.575 123.390 142.275 124.790 ;
        RECT 142.575 123.390 144.275 124.790 ;
        RECT 144.575 123.390 146.275 124.790 ;
        RECT 146.575 123.390 148.275 124.790 ;
        RECT 148.575 123.390 150.275 124.790 ;
        RECT 150.575 123.390 152.275 124.790 ;
        RECT 152.575 123.390 154.275 124.790 ;
        RECT 6.840 121.540 8.540 122.940 ;
        RECT 8.840 121.540 10.540 122.940 ;
        RECT 10.840 121.540 12.540 122.940 ;
        RECT 12.840 121.540 14.540 122.940 ;
        RECT 14.840 121.540 16.540 122.940 ;
        RECT 16.840 121.540 18.540 122.940 ;
        RECT 18.840 121.540 20.540 122.940 ;
        RECT 20.840 121.540 22.540 122.940 ;
        RECT 22.840 121.540 24.540 122.940 ;
        RECT 24.840 121.540 26.540 122.940 ;
        RECT 26.840 121.540 28.540 122.940 ;
        RECT 28.840 121.540 30.540 122.940 ;
        RECT 30.840 121.540 32.540 122.940 ;
        RECT 32.840 121.540 34.540 122.940 ;
        RECT 34.840 121.540 36.540 122.940 ;
        RECT 36.840 121.540 38.540 122.940 ;
        RECT 38.840 121.540 40.540 122.940 ;
        RECT 40.840 121.540 42.540 122.940 ;
        RECT 42.840 121.540 44.540 122.940 ;
        RECT 44.840 121.540 46.540 122.940 ;
        RECT 46.840 121.540 48.540 122.940 ;
        RECT 48.840 121.540 50.540 122.940 ;
        RECT 50.840 121.540 52.540 122.940 ;
        RECT 52.840 121.540 54.540 122.940 ;
        RECT 54.840 121.540 56.540 122.940 ;
        RECT 56.840 121.540 58.540 122.940 ;
        RECT 58.840 121.540 60.540 122.940 ;
        RECT 60.840 121.540 62.540 122.940 ;
        RECT 62.840 121.540 64.540 122.940 ;
        RECT 64.840 121.540 66.540 122.940 ;
        RECT 66.840 121.540 68.540 122.940 ;
        RECT 68.840 121.540 70.540 122.940 ;
        RECT 70.840 121.540 72.540 122.940 ;
        RECT 72.840 121.540 74.540 122.940 ;
        RECT 86.575 121.540 88.275 122.940 ;
        RECT 88.575 121.540 90.275 122.940 ;
        RECT 90.575 121.540 92.275 122.940 ;
        RECT 92.575 121.540 94.275 122.940 ;
        RECT 94.575 121.540 96.275 122.940 ;
        RECT 96.575 121.540 98.275 122.940 ;
        RECT 98.575 121.540 100.275 122.940 ;
        RECT 100.575 121.540 102.275 122.940 ;
        RECT 102.575 121.540 104.275 122.940 ;
        RECT 104.575 121.540 106.275 122.940 ;
        RECT 106.575 121.540 108.275 122.940 ;
        RECT 108.575 121.540 110.275 122.940 ;
        RECT 110.575 121.540 112.275 122.940 ;
        RECT 112.575 121.540 114.275 122.940 ;
        RECT 114.575 121.540 116.275 122.940 ;
        RECT 116.575 121.540 118.275 122.940 ;
        RECT 118.575 121.540 120.275 122.940 ;
        RECT 120.575 121.540 122.275 122.940 ;
        RECT 122.575 121.540 124.275 122.940 ;
        RECT 124.575 121.540 126.275 122.940 ;
        RECT 126.575 121.540 128.275 122.940 ;
        RECT 128.575 121.540 130.275 122.940 ;
        RECT 130.575 121.540 132.275 122.940 ;
        RECT 132.575 121.540 134.275 122.940 ;
        RECT 134.575 121.540 136.275 122.940 ;
        RECT 136.575 121.540 138.275 122.940 ;
        RECT 138.575 121.540 140.275 122.940 ;
        RECT 140.575 121.540 142.275 122.940 ;
        RECT 142.575 121.540 144.275 122.940 ;
        RECT 144.575 121.540 146.275 122.940 ;
        RECT 146.575 121.540 148.275 122.940 ;
        RECT 148.575 121.540 150.275 122.940 ;
        RECT 150.575 121.540 152.275 122.940 ;
        RECT 152.575 121.540 154.275 122.940 ;
        RECT 6.840 119.690 8.540 121.090 ;
        RECT 8.840 119.690 10.540 121.090 ;
        RECT 10.840 119.690 12.540 121.090 ;
        RECT 12.840 119.690 14.540 121.090 ;
        RECT 14.840 119.690 16.540 121.090 ;
        RECT 16.840 119.690 18.540 121.090 ;
        RECT 18.840 119.690 20.540 121.090 ;
        RECT 20.840 119.690 22.540 121.090 ;
        RECT 22.840 119.690 24.540 121.090 ;
        RECT 24.840 119.690 26.540 121.090 ;
        RECT 26.840 119.690 28.540 121.090 ;
        RECT 28.840 119.690 30.540 121.090 ;
        RECT 30.840 119.690 32.540 121.090 ;
        RECT 32.840 119.690 34.540 121.090 ;
        RECT 34.840 119.690 36.540 121.090 ;
        RECT 36.840 119.690 38.540 121.090 ;
        RECT 38.840 119.690 40.540 121.090 ;
        RECT 40.840 119.690 42.540 121.090 ;
        RECT 42.840 119.690 44.540 121.090 ;
        RECT 44.840 119.690 46.540 121.090 ;
        RECT 46.840 119.690 48.540 121.090 ;
        RECT 48.840 119.690 50.540 121.090 ;
        RECT 50.840 119.690 52.540 121.090 ;
        RECT 52.840 119.690 54.540 121.090 ;
        RECT 54.840 119.690 56.540 121.090 ;
        RECT 56.840 119.690 58.540 121.090 ;
        RECT 58.840 119.690 60.540 121.090 ;
        RECT 60.840 119.690 62.540 121.090 ;
        RECT 62.840 119.690 64.540 121.090 ;
        RECT 64.840 119.690 66.540 121.090 ;
        RECT 66.840 119.690 68.540 121.090 ;
        RECT 68.840 119.690 70.540 121.090 ;
        RECT 70.840 119.690 72.540 121.090 ;
        RECT 72.840 119.690 74.540 121.090 ;
        RECT 86.575 119.690 88.275 121.090 ;
        RECT 88.575 119.690 90.275 121.090 ;
        RECT 90.575 119.690 92.275 121.090 ;
        RECT 92.575 119.690 94.275 121.090 ;
        RECT 94.575 119.690 96.275 121.090 ;
        RECT 96.575 119.690 98.275 121.090 ;
        RECT 98.575 119.690 100.275 121.090 ;
        RECT 100.575 119.690 102.275 121.090 ;
        RECT 102.575 119.690 104.275 121.090 ;
        RECT 104.575 119.690 106.275 121.090 ;
        RECT 106.575 119.690 108.275 121.090 ;
        RECT 108.575 119.690 110.275 121.090 ;
        RECT 110.575 119.690 112.275 121.090 ;
        RECT 112.575 119.690 114.275 121.090 ;
        RECT 114.575 119.690 116.275 121.090 ;
        RECT 116.575 119.690 118.275 121.090 ;
        RECT 118.575 119.690 120.275 121.090 ;
        RECT 120.575 119.690 122.275 121.090 ;
        RECT 122.575 119.690 124.275 121.090 ;
        RECT 124.575 119.690 126.275 121.090 ;
        RECT 126.575 119.690 128.275 121.090 ;
        RECT 128.575 119.690 130.275 121.090 ;
        RECT 130.575 119.690 132.275 121.090 ;
        RECT 132.575 119.690 134.275 121.090 ;
        RECT 134.575 119.690 136.275 121.090 ;
        RECT 136.575 119.690 138.275 121.090 ;
        RECT 138.575 119.690 140.275 121.090 ;
        RECT 140.575 119.690 142.275 121.090 ;
        RECT 142.575 119.690 144.275 121.090 ;
        RECT 144.575 119.690 146.275 121.090 ;
        RECT 146.575 119.690 148.275 121.090 ;
        RECT 148.575 119.690 150.275 121.090 ;
        RECT 150.575 119.690 152.275 121.090 ;
        RECT 152.575 119.690 154.275 121.090 ;
        RECT 6.840 117.840 8.540 119.240 ;
        RECT 8.840 117.840 10.540 119.240 ;
        RECT 10.840 117.840 12.540 119.240 ;
        RECT 12.840 117.840 14.540 119.240 ;
        RECT 14.840 117.840 16.540 119.240 ;
        RECT 16.840 117.840 18.540 119.240 ;
        RECT 18.840 117.840 20.540 119.240 ;
        RECT 20.840 117.840 22.540 119.240 ;
        RECT 22.840 117.840 24.540 119.240 ;
        RECT 24.840 117.840 26.540 119.240 ;
        RECT 26.840 117.840 28.540 119.240 ;
        RECT 28.840 117.840 30.540 119.240 ;
        RECT 30.840 117.840 32.540 119.240 ;
        RECT 32.840 117.840 34.540 119.240 ;
        RECT 34.840 117.840 36.540 119.240 ;
        RECT 36.840 117.840 38.540 119.240 ;
        RECT 38.840 117.840 40.540 119.240 ;
        RECT 40.840 117.840 42.540 119.240 ;
        RECT 42.840 117.840 44.540 119.240 ;
        RECT 44.840 117.840 46.540 119.240 ;
        RECT 46.840 117.840 48.540 119.240 ;
        RECT 48.840 117.840 50.540 119.240 ;
        RECT 50.840 117.840 52.540 119.240 ;
        RECT 52.840 117.840 54.540 119.240 ;
        RECT 54.840 117.840 56.540 119.240 ;
        RECT 56.840 117.840 58.540 119.240 ;
        RECT 58.840 117.840 60.540 119.240 ;
        RECT 60.840 117.840 62.540 119.240 ;
        RECT 62.840 117.840 64.540 119.240 ;
        RECT 64.840 117.840 66.540 119.240 ;
        RECT 66.840 117.840 68.540 119.240 ;
        RECT 68.840 117.840 70.540 119.240 ;
        RECT 70.840 117.840 72.540 119.240 ;
        RECT 72.840 117.840 74.540 119.240 ;
        RECT 86.575 117.840 88.275 119.240 ;
        RECT 88.575 117.840 90.275 119.240 ;
        RECT 90.575 117.840 92.275 119.240 ;
        RECT 92.575 117.840 94.275 119.240 ;
        RECT 94.575 117.840 96.275 119.240 ;
        RECT 96.575 117.840 98.275 119.240 ;
        RECT 98.575 117.840 100.275 119.240 ;
        RECT 100.575 117.840 102.275 119.240 ;
        RECT 102.575 117.840 104.275 119.240 ;
        RECT 104.575 117.840 106.275 119.240 ;
        RECT 106.575 117.840 108.275 119.240 ;
        RECT 108.575 117.840 110.275 119.240 ;
        RECT 110.575 117.840 112.275 119.240 ;
        RECT 112.575 117.840 114.275 119.240 ;
        RECT 114.575 117.840 116.275 119.240 ;
        RECT 116.575 117.840 118.275 119.240 ;
        RECT 118.575 117.840 120.275 119.240 ;
        RECT 120.575 117.840 122.275 119.240 ;
        RECT 122.575 117.840 124.275 119.240 ;
        RECT 124.575 117.840 126.275 119.240 ;
        RECT 126.575 117.840 128.275 119.240 ;
        RECT 128.575 117.840 130.275 119.240 ;
        RECT 130.575 117.840 132.275 119.240 ;
        RECT 132.575 117.840 134.275 119.240 ;
        RECT 134.575 117.840 136.275 119.240 ;
        RECT 136.575 117.840 138.275 119.240 ;
        RECT 138.575 117.840 140.275 119.240 ;
        RECT 140.575 117.840 142.275 119.240 ;
        RECT 142.575 117.840 144.275 119.240 ;
        RECT 144.575 117.840 146.275 119.240 ;
        RECT 146.575 117.840 148.275 119.240 ;
        RECT 148.575 117.840 150.275 119.240 ;
        RECT 150.575 117.840 152.275 119.240 ;
        RECT 152.575 117.840 154.275 119.240 ;
        RECT 6.840 115.990 8.540 117.390 ;
        RECT 8.840 115.990 10.540 117.390 ;
        RECT 10.840 115.990 12.540 117.390 ;
        RECT 12.840 115.990 14.540 117.390 ;
        RECT 14.840 115.990 16.540 117.390 ;
        RECT 16.840 115.990 18.540 117.390 ;
        RECT 18.840 115.990 20.540 117.390 ;
        RECT 20.840 115.990 22.540 117.390 ;
        RECT 22.840 115.990 24.540 117.390 ;
        RECT 24.840 115.990 26.540 117.390 ;
        RECT 26.840 115.990 28.540 117.390 ;
        RECT 28.840 115.990 30.540 117.390 ;
        RECT 30.840 115.990 32.540 117.390 ;
        RECT 32.840 115.990 34.540 117.390 ;
        RECT 34.840 115.990 36.540 117.390 ;
        RECT 36.840 115.990 38.540 117.390 ;
        RECT 38.840 115.990 40.540 117.390 ;
        RECT 40.840 115.990 42.540 117.390 ;
        RECT 42.840 115.990 44.540 117.390 ;
        RECT 44.840 115.990 46.540 117.390 ;
        RECT 46.840 115.990 48.540 117.390 ;
        RECT 48.840 115.990 50.540 117.390 ;
        RECT 50.840 115.990 52.540 117.390 ;
        RECT 52.840 115.990 54.540 117.390 ;
        RECT 54.840 115.990 56.540 117.390 ;
        RECT 56.840 115.990 58.540 117.390 ;
        RECT 58.840 115.990 60.540 117.390 ;
        RECT 60.840 115.990 62.540 117.390 ;
        RECT 62.840 115.990 64.540 117.390 ;
        RECT 64.840 115.990 66.540 117.390 ;
        RECT 66.840 115.990 68.540 117.390 ;
        RECT 68.840 115.990 70.540 117.390 ;
        RECT 70.840 115.990 72.540 117.390 ;
        RECT 72.840 115.990 74.540 117.390 ;
        RECT 86.575 115.990 88.275 117.390 ;
        RECT 88.575 115.990 90.275 117.390 ;
        RECT 90.575 115.990 92.275 117.390 ;
        RECT 92.575 115.990 94.275 117.390 ;
        RECT 94.575 115.990 96.275 117.390 ;
        RECT 96.575 115.990 98.275 117.390 ;
        RECT 98.575 115.990 100.275 117.390 ;
        RECT 100.575 115.990 102.275 117.390 ;
        RECT 102.575 115.990 104.275 117.390 ;
        RECT 104.575 115.990 106.275 117.390 ;
        RECT 106.575 115.990 108.275 117.390 ;
        RECT 108.575 115.990 110.275 117.390 ;
        RECT 110.575 115.990 112.275 117.390 ;
        RECT 112.575 115.990 114.275 117.390 ;
        RECT 114.575 115.990 116.275 117.390 ;
        RECT 116.575 115.990 118.275 117.390 ;
        RECT 118.575 115.990 120.275 117.390 ;
        RECT 120.575 115.990 122.275 117.390 ;
        RECT 122.575 115.990 124.275 117.390 ;
        RECT 124.575 115.990 126.275 117.390 ;
        RECT 126.575 115.990 128.275 117.390 ;
        RECT 128.575 115.990 130.275 117.390 ;
        RECT 130.575 115.990 132.275 117.390 ;
        RECT 132.575 115.990 134.275 117.390 ;
        RECT 134.575 115.990 136.275 117.390 ;
        RECT 136.575 115.990 138.275 117.390 ;
        RECT 138.575 115.990 140.275 117.390 ;
        RECT 140.575 115.990 142.275 117.390 ;
        RECT 142.575 115.990 144.275 117.390 ;
        RECT 144.575 115.990 146.275 117.390 ;
        RECT 146.575 115.990 148.275 117.390 ;
        RECT 148.575 115.990 150.275 117.390 ;
        RECT 150.575 115.990 152.275 117.390 ;
        RECT 152.575 115.990 154.275 117.390 ;
        RECT 6.840 114.140 8.540 115.540 ;
        RECT 8.840 114.140 10.540 115.540 ;
        RECT 10.840 114.140 12.540 115.540 ;
        RECT 12.840 114.140 14.540 115.540 ;
        RECT 14.840 114.140 16.540 115.540 ;
        RECT 16.840 114.140 18.540 115.540 ;
        RECT 18.840 114.140 20.540 115.540 ;
        RECT 20.840 114.140 22.540 115.540 ;
        RECT 22.840 114.140 24.540 115.540 ;
        RECT 24.840 114.140 26.540 115.540 ;
        RECT 26.840 114.140 28.540 115.540 ;
        RECT 28.840 114.140 30.540 115.540 ;
        RECT 30.840 114.140 32.540 115.540 ;
        RECT 32.840 114.140 34.540 115.540 ;
        RECT 34.840 114.140 36.540 115.540 ;
        RECT 36.840 114.140 38.540 115.540 ;
        RECT 38.840 114.140 40.540 115.540 ;
        RECT 40.840 114.140 42.540 115.540 ;
        RECT 42.840 114.140 44.540 115.540 ;
        RECT 44.840 114.140 46.540 115.540 ;
        RECT 46.840 114.140 48.540 115.540 ;
        RECT 48.840 114.140 50.540 115.540 ;
        RECT 50.840 114.140 52.540 115.540 ;
        RECT 52.840 114.140 54.540 115.540 ;
        RECT 54.840 114.140 56.540 115.540 ;
        RECT 56.840 114.140 58.540 115.540 ;
        RECT 58.840 114.140 60.540 115.540 ;
        RECT 60.840 114.140 62.540 115.540 ;
        RECT 62.840 114.140 64.540 115.540 ;
        RECT 64.840 114.140 66.540 115.540 ;
        RECT 66.840 114.140 68.540 115.540 ;
        RECT 68.840 114.140 70.540 115.540 ;
        RECT 70.840 114.140 72.540 115.540 ;
        RECT 72.840 114.140 74.540 115.540 ;
        RECT 86.575 114.140 88.275 115.540 ;
        RECT 88.575 114.140 90.275 115.540 ;
        RECT 90.575 114.140 92.275 115.540 ;
        RECT 92.575 114.140 94.275 115.540 ;
        RECT 94.575 114.140 96.275 115.540 ;
        RECT 96.575 114.140 98.275 115.540 ;
        RECT 98.575 114.140 100.275 115.540 ;
        RECT 100.575 114.140 102.275 115.540 ;
        RECT 102.575 114.140 104.275 115.540 ;
        RECT 104.575 114.140 106.275 115.540 ;
        RECT 106.575 114.140 108.275 115.540 ;
        RECT 108.575 114.140 110.275 115.540 ;
        RECT 110.575 114.140 112.275 115.540 ;
        RECT 112.575 114.140 114.275 115.540 ;
        RECT 114.575 114.140 116.275 115.540 ;
        RECT 116.575 114.140 118.275 115.540 ;
        RECT 118.575 114.140 120.275 115.540 ;
        RECT 120.575 114.140 122.275 115.540 ;
        RECT 122.575 114.140 124.275 115.540 ;
        RECT 124.575 114.140 126.275 115.540 ;
        RECT 126.575 114.140 128.275 115.540 ;
        RECT 128.575 114.140 130.275 115.540 ;
        RECT 130.575 114.140 132.275 115.540 ;
        RECT 132.575 114.140 134.275 115.540 ;
        RECT 134.575 114.140 136.275 115.540 ;
        RECT 136.575 114.140 138.275 115.540 ;
        RECT 138.575 114.140 140.275 115.540 ;
        RECT 140.575 114.140 142.275 115.540 ;
        RECT 142.575 114.140 144.275 115.540 ;
        RECT 144.575 114.140 146.275 115.540 ;
        RECT 146.575 114.140 148.275 115.540 ;
        RECT 148.575 114.140 150.275 115.540 ;
        RECT 150.575 114.140 152.275 115.540 ;
        RECT 152.575 114.140 154.275 115.540 ;
        RECT 6.840 112.290 8.540 113.690 ;
        RECT 8.840 112.290 10.540 113.690 ;
        RECT 10.840 112.290 12.540 113.690 ;
        RECT 12.840 112.290 14.540 113.690 ;
        RECT 14.840 112.290 16.540 113.690 ;
        RECT 16.840 112.290 18.540 113.690 ;
        RECT 18.840 112.290 20.540 113.690 ;
        RECT 20.840 112.290 22.540 113.690 ;
        RECT 22.840 112.290 24.540 113.690 ;
        RECT 24.840 112.290 26.540 113.690 ;
        RECT 26.840 112.290 28.540 113.690 ;
        RECT 28.840 112.290 30.540 113.690 ;
        RECT 30.840 112.290 32.540 113.690 ;
        RECT 32.840 112.290 34.540 113.690 ;
        RECT 34.840 112.290 36.540 113.690 ;
        RECT 36.840 112.290 38.540 113.690 ;
        RECT 38.840 112.290 40.540 113.690 ;
        RECT 40.840 112.290 42.540 113.690 ;
        RECT 42.840 112.290 44.540 113.690 ;
        RECT 44.840 112.290 46.540 113.690 ;
        RECT 46.840 112.290 48.540 113.690 ;
        RECT 48.840 112.290 50.540 113.690 ;
        RECT 50.840 112.290 52.540 113.690 ;
        RECT 52.840 112.290 54.540 113.690 ;
        RECT 54.840 112.290 56.540 113.690 ;
        RECT 56.840 112.290 58.540 113.690 ;
        RECT 58.840 112.290 60.540 113.690 ;
        RECT 60.840 112.290 62.540 113.690 ;
        RECT 62.840 112.290 64.540 113.690 ;
        RECT 64.840 112.290 66.540 113.690 ;
        RECT 66.840 112.290 68.540 113.690 ;
        RECT 68.840 112.290 70.540 113.690 ;
        RECT 70.840 112.290 72.540 113.690 ;
        RECT 72.840 112.290 74.540 113.690 ;
        RECT 86.575 112.290 88.275 113.690 ;
        RECT 88.575 112.290 90.275 113.690 ;
        RECT 90.575 112.290 92.275 113.690 ;
        RECT 92.575 112.290 94.275 113.690 ;
        RECT 94.575 112.290 96.275 113.690 ;
        RECT 96.575 112.290 98.275 113.690 ;
        RECT 98.575 112.290 100.275 113.690 ;
        RECT 100.575 112.290 102.275 113.690 ;
        RECT 102.575 112.290 104.275 113.690 ;
        RECT 104.575 112.290 106.275 113.690 ;
        RECT 106.575 112.290 108.275 113.690 ;
        RECT 108.575 112.290 110.275 113.690 ;
        RECT 110.575 112.290 112.275 113.690 ;
        RECT 112.575 112.290 114.275 113.690 ;
        RECT 114.575 112.290 116.275 113.690 ;
        RECT 116.575 112.290 118.275 113.690 ;
        RECT 118.575 112.290 120.275 113.690 ;
        RECT 120.575 112.290 122.275 113.690 ;
        RECT 122.575 112.290 124.275 113.690 ;
        RECT 124.575 112.290 126.275 113.690 ;
        RECT 126.575 112.290 128.275 113.690 ;
        RECT 128.575 112.290 130.275 113.690 ;
        RECT 130.575 112.290 132.275 113.690 ;
        RECT 132.575 112.290 134.275 113.690 ;
        RECT 134.575 112.290 136.275 113.690 ;
        RECT 136.575 112.290 138.275 113.690 ;
        RECT 138.575 112.290 140.275 113.690 ;
        RECT 140.575 112.290 142.275 113.690 ;
        RECT 142.575 112.290 144.275 113.690 ;
        RECT 144.575 112.290 146.275 113.690 ;
        RECT 146.575 112.290 148.275 113.690 ;
        RECT 148.575 112.290 150.275 113.690 ;
        RECT 150.575 112.290 152.275 113.690 ;
        RECT 152.575 112.290 154.275 113.690 ;
        RECT 6.840 110.440 8.540 111.840 ;
        RECT 8.840 110.440 10.540 111.840 ;
        RECT 10.840 110.440 12.540 111.840 ;
        RECT 12.840 110.440 14.540 111.840 ;
        RECT 14.840 110.440 16.540 111.840 ;
        RECT 16.840 110.440 18.540 111.840 ;
        RECT 18.840 110.440 20.540 111.840 ;
        RECT 20.840 110.440 22.540 111.840 ;
        RECT 22.840 110.440 24.540 111.840 ;
        RECT 24.840 110.440 26.540 111.840 ;
        RECT 26.840 110.440 28.540 111.840 ;
        RECT 28.840 110.440 30.540 111.840 ;
        RECT 30.840 110.440 32.540 111.840 ;
        RECT 32.840 110.440 34.540 111.840 ;
        RECT 34.840 110.440 36.540 111.840 ;
        RECT 36.840 110.440 38.540 111.840 ;
        RECT 38.840 110.440 40.540 111.840 ;
        RECT 40.840 110.440 42.540 111.840 ;
        RECT 42.840 110.440 44.540 111.840 ;
        RECT 44.840 110.440 46.540 111.840 ;
        RECT 46.840 110.440 48.540 111.840 ;
        RECT 48.840 110.440 50.540 111.840 ;
        RECT 50.840 110.440 52.540 111.840 ;
        RECT 52.840 110.440 54.540 111.840 ;
        RECT 54.840 110.440 56.540 111.840 ;
        RECT 56.840 110.440 58.540 111.840 ;
        RECT 58.840 110.440 60.540 111.840 ;
        RECT 60.840 110.440 62.540 111.840 ;
        RECT 62.840 110.440 64.540 111.840 ;
        RECT 64.840 110.440 66.540 111.840 ;
        RECT 66.840 110.440 68.540 111.840 ;
        RECT 68.840 110.440 70.540 111.840 ;
        RECT 70.840 110.440 72.540 111.840 ;
        RECT 72.840 110.440 74.540 111.840 ;
        RECT 86.575 110.440 88.275 111.840 ;
        RECT 88.575 110.440 90.275 111.840 ;
        RECT 90.575 110.440 92.275 111.840 ;
        RECT 92.575 110.440 94.275 111.840 ;
        RECT 94.575 110.440 96.275 111.840 ;
        RECT 96.575 110.440 98.275 111.840 ;
        RECT 98.575 110.440 100.275 111.840 ;
        RECT 100.575 110.440 102.275 111.840 ;
        RECT 102.575 110.440 104.275 111.840 ;
        RECT 104.575 110.440 106.275 111.840 ;
        RECT 106.575 110.440 108.275 111.840 ;
        RECT 108.575 110.440 110.275 111.840 ;
        RECT 110.575 110.440 112.275 111.840 ;
        RECT 112.575 110.440 114.275 111.840 ;
        RECT 114.575 110.440 116.275 111.840 ;
        RECT 116.575 110.440 118.275 111.840 ;
        RECT 118.575 110.440 120.275 111.840 ;
        RECT 120.575 110.440 122.275 111.840 ;
        RECT 122.575 110.440 124.275 111.840 ;
        RECT 124.575 110.440 126.275 111.840 ;
        RECT 126.575 110.440 128.275 111.840 ;
        RECT 128.575 110.440 130.275 111.840 ;
        RECT 130.575 110.440 132.275 111.840 ;
        RECT 132.575 110.440 134.275 111.840 ;
        RECT 134.575 110.440 136.275 111.840 ;
        RECT 136.575 110.440 138.275 111.840 ;
        RECT 138.575 110.440 140.275 111.840 ;
        RECT 140.575 110.440 142.275 111.840 ;
        RECT 142.575 110.440 144.275 111.840 ;
        RECT 144.575 110.440 146.275 111.840 ;
        RECT 146.575 110.440 148.275 111.840 ;
        RECT 148.575 110.440 150.275 111.840 ;
        RECT 150.575 110.440 152.275 111.840 ;
        RECT 152.575 110.440 154.275 111.840 ;
        RECT 6.840 108.590 8.540 109.990 ;
        RECT 8.840 108.590 10.540 109.990 ;
        RECT 10.840 108.590 12.540 109.990 ;
        RECT 12.840 108.590 14.540 109.990 ;
        RECT 14.840 108.590 16.540 109.990 ;
        RECT 16.840 108.590 18.540 109.990 ;
        RECT 18.840 108.590 20.540 109.990 ;
        RECT 20.840 108.590 22.540 109.990 ;
        RECT 22.840 108.590 24.540 109.990 ;
        RECT 24.840 108.590 26.540 109.990 ;
        RECT 26.840 108.590 28.540 109.990 ;
        RECT 28.840 108.590 30.540 109.990 ;
        RECT 30.840 108.590 32.540 109.990 ;
        RECT 32.840 108.590 34.540 109.990 ;
        RECT 34.840 108.590 36.540 109.990 ;
        RECT 36.840 108.590 38.540 109.990 ;
        RECT 38.840 108.590 40.540 109.990 ;
        RECT 40.840 108.590 42.540 109.990 ;
        RECT 42.840 108.590 44.540 109.990 ;
        RECT 44.840 108.590 46.540 109.990 ;
        RECT 46.840 108.590 48.540 109.990 ;
        RECT 48.840 108.590 50.540 109.990 ;
        RECT 50.840 108.590 52.540 109.990 ;
        RECT 52.840 108.590 54.540 109.990 ;
        RECT 54.840 108.590 56.540 109.990 ;
        RECT 56.840 108.590 58.540 109.990 ;
        RECT 58.840 108.590 60.540 109.990 ;
        RECT 60.840 108.590 62.540 109.990 ;
        RECT 62.840 108.590 64.540 109.990 ;
        RECT 64.840 108.590 66.540 109.990 ;
        RECT 66.840 108.590 68.540 109.990 ;
        RECT 68.840 108.590 70.540 109.990 ;
        RECT 70.840 108.590 72.540 109.990 ;
        RECT 72.840 108.590 74.540 109.990 ;
        RECT 86.575 108.590 88.275 109.990 ;
        RECT 88.575 108.590 90.275 109.990 ;
        RECT 90.575 108.590 92.275 109.990 ;
        RECT 92.575 108.590 94.275 109.990 ;
        RECT 94.575 108.590 96.275 109.990 ;
        RECT 96.575 108.590 98.275 109.990 ;
        RECT 98.575 108.590 100.275 109.990 ;
        RECT 100.575 108.590 102.275 109.990 ;
        RECT 102.575 108.590 104.275 109.990 ;
        RECT 104.575 108.590 106.275 109.990 ;
        RECT 106.575 108.590 108.275 109.990 ;
        RECT 108.575 108.590 110.275 109.990 ;
        RECT 110.575 108.590 112.275 109.990 ;
        RECT 112.575 108.590 114.275 109.990 ;
        RECT 114.575 108.590 116.275 109.990 ;
        RECT 116.575 108.590 118.275 109.990 ;
        RECT 118.575 108.590 120.275 109.990 ;
        RECT 120.575 108.590 122.275 109.990 ;
        RECT 122.575 108.590 124.275 109.990 ;
        RECT 124.575 108.590 126.275 109.990 ;
        RECT 126.575 108.590 128.275 109.990 ;
        RECT 128.575 108.590 130.275 109.990 ;
        RECT 130.575 108.590 132.275 109.990 ;
        RECT 132.575 108.590 134.275 109.990 ;
        RECT 134.575 108.590 136.275 109.990 ;
        RECT 136.575 108.590 138.275 109.990 ;
        RECT 138.575 108.590 140.275 109.990 ;
        RECT 140.575 108.590 142.275 109.990 ;
        RECT 142.575 108.590 144.275 109.990 ;
        RECT 144.575 108.590 146.275 109.990 ;
        RECT 146.575 108.590 148.275 109.990 ;
        RECT 148.575 108.590 150.275 109.990 ;
        RECT 150.575 108.590 152.275 109.990 ;
        RECT 152.575 108.590 154.275 109.990 ;
        RECT 6.840 106.740 8.540 108.140 ;
        RECT 8.840 106.740 10.540 108.140 ;
        RECT 10.840 106.740 12.540 108.140 ;
        RECT 12.840 106.740 14.540 108.140 ;
        RECT 14.840 106.740 16.540 108.140 ;
        RECT 16.840 106.740 18.540 108.140 ;
        RECT 18.840 106.740 20.540 108.140 ;
        RECT 20.840 106.740 22.540 108.140 ;
        RECT 22.840 106.740 24.540 108.140 ;
        RECT 24.840 106.740 26.540 108.140 ;
        RECT 26.840 106.740 28.540 108.140 ;
        RECT 28.840 106.740 30.540 108.140 ;
        RECT 30.840 106.740 32.540 108.140 ;
        RECT 32.840 106.740 34.540 108.140 ;
        RECT 34.840 106.740 36.540 108.140 ;
        RECT 36.840 106.740 38.540 108.140 ;
        RECT 38.840 106.740 40.540 108.140 ;
        RECT 40.840 106.740 42.540 108.140 ;
        RECT 42.840 106.740 44.540 108.140 ;
        RECT 44.840 106.740 46.540 108.140 ;
        RECT 46.840 106.740 48.540 108.140 ;
        RECT 48.840 106.740 50.540 108.140 ;
        RECT 50.840 106.740 52.540 108.140 ;
        RECT 52.840 106.740 54.540 108.140 ;
        RECT 54.840 106.740 56.540 108.140 ;
        RECT 56.840 106.740 58.540 108.140 ;
        RECT 58.840 106.740 60.540 108.140 ;
        RECT 60.840 106.740 62.540 108.140 ;
        RECT 62.840 106.740 64.540 108.140 ;
        RECT 64.840 106.740 66.540 108.140 ;
        RECT 66.840 106.740 68.540 108.140 ;
        RECT 68.840 106.740 70.540 108.140 ;
        RECT 70.840 106.740 72.540 108.140 ;
        RECT 72.840 106.740 74.540 108.140 ;
        RECT 86.575 106.740 88.275 108.140 ;
        RECT 88.575 106.740 90.275 108.140 ;
        RECT 90.575 106.740 92.275 108.140 ;
        RECT 92.575 106.740 94.275 108.140 ;
        RECT 94.575 106.740 96.275 108.140 ;
        RECT 96.575 106.740 98.275 108.140 ;
        RECT 98.575 106.740 100.275 108.140 ;
        RECT 100.575 106.740 102.275 108.140 ;
        RECT 102.575 106.740 104.275 108.140 ;
        RECT 104.575 106.740 106.275 108.140 ;
        RECT 106.575 106.740 108.275 108.140 ;
        RECT 108.575 106.740 110.275 108.140 ;
        RECT 110.575 106.740 112.275 108.140 ;
        RECT 112.575 106.740 114.275 108.140 ;
        RECT 114.575 106.740 116.275 108.140 ;
        RECT 116.575 106.740 118.275 108.140 ;
        RECT 118.575 106.740 120.275 108.140 ;
        RECT 120.575 106.740 122.275 108.140 ;
        RECT 122.575 106.740 124.275 108.140 ;
        RECT 124.575 106.740 126.275 108.140 ;
        RECT 126.575 106.740 128.275 108.140 ;
        RECT 128.575 106.740 130.275 108.140 ;
        RECT 130.575 106.740 132.275 108.140 ;
        RECT 132.575 106.740 134.275 108.140 ;
        RECT 134.575 106.740 136.275 108.140 ;
        RECT 136.575 106.740 138.275 108.140 ;
        RECT 138.575 106.740 140.275 108.140 ;
        RECT 140.575 106.740 142.275 108.140 ;
        RECT 142.575 106.740 144.275 108.140 ;
        RECT 144.575 106.740 146.275 108.140 ;
        RECT 146.575 106.740 148.275 108.140 ;
        RECT 148.575 106.740 150.275 108.140 ;
        RECT 150.575 106.740 152.275 108.140 ;
        RECT 152.575 106.740 154.275 108.140 ;
        RECT 6.840 104.890 8.540 106.290 ;
        RECT 8.840 104.890 10.540 106.290 ;
        RECT 10.840 104.890 12.540 106.290 ;
        RECT 12.840 104.890 14.540 106.290 ;
        RECT 14.840 104.890 16.540 106.290 ;
        RECT 16.840 104.890 18.540 106.290 ;
        RECT 18.840 104.890 20.540 106.290 ;
        RECT 20.840 104.890 22.540 106.290 ;
        RECT 22.840 104.890 24.540 106.290 ;
        RECT 24.840 104.890 26.540 106.290 ;
        RECT 26.840 104.890 28.540 106.290 ;
        RECT 28.840 104.890 30.540 106.290 ;
        RECT 30.840 104.890 32.540 106.290 ;
        RECT 32.840 104.890 34.540 106.290 ;
        RECT 34.840 104.890 36.540 106.290 ;
        RECT 36.840 104.890 38.540 106.290 ;
        RECT 38.840 104.890 40.540 106.290 ;
        RECT 40.840 104.890 42.540 106.290 ;
        RECT 42.840 104.890 44.540 106.290 ;
        RECT 44.840 104.890 46.540 106.290 ;
        RECT 46.840 104.890 48.540 106.290 ;
        RECT 48.840 104.890 50.540 106.290 ;
        RECT 50.840 104.890 52.540 106.290 ;
        RECT 52.840 104.890 54.540 106.290 ;
        RECT 54.840 104.890 56.540 106.290 ;
        RECT 56.840 104.890 58.540 106.290 ;
        RECT 58.840 104.890 60.540 106.290 ;
        RECT 60.840 104.890 62.540 106.290 ;
        RECT 62.840 104.890 64.540 106.290 ;
        RECT 64.840 104.890 66.540 106.290 ;
        RECT 66.840 104.890 68.540 106.290 ;
        RECT 68.840 104.890 70.540 106.290 ;
        RECT 70.840 104.890 72.540 106.290 ;
        RECT 72.840 104.890 74.540 106.290 ;
        RECT 86.575 104.890 88.275 106.290 ;
        RECT 88.575 104.890 90.275 106.290 ;
        RECT 90.575 104.890 92.275 106.290 ;
        RECT 92.575 104.890 94.275 106.290 ;
        RECT 94.575 104.890 96.275 106.290 ;
        RECT 96.575 104.890 98.275 106.290 ;
        RECT 98.575 104.890 100.275 106.290 ;
        RECT 100.575 104.890 102.275 106.290 ;
        RECT 102.575 104.890 104.275 106.290 ;
        RECT 104.575 104.890 106.275 106.290 ;
        RECT 106.575 104.890 108.275 106.290 ;
        RECT 108.575 104.890 110.275 106.290 ;
        RECT 110.575 104.890 112.275 106.290 ;
        RECT 112.575 104.890 114.275 106.290 ;
        RECT 114.575 104.890 116.275 106.290 ;
        RECT 116.575 104.890 118.275 106.290 ;
        RECT 118.575 104.890 120.275 106.290 ;
        RECT 120.575 104.890 122.275 106.290 ;
        RECT 122.575 104.890 124.275 106.290 ;
        RECT 124.575 104.890 126.275 106.290 ;
        RECT 126.575 104.890 128.275 106.290 ;
        RECT 128.575 104.890 130.275 106.290 ;
        RECT 130.575 104.890 132.275 106.290 ;
        RECT 132.575 104.890 134.275 106.290 ;
        RECT 134.575 104.890 136.275 106.290 ;
        RECT 136.575 104.890 138.275 106.290 ;
        RECT 138.575 104.890 140.275 106.290 ;
        RECT 140.575 104.890 142.275 106.290 ;
        RECT 142.575 104.890 144.275 106.290 ;
        RECT 144.575 104.890 146.275 106.290 ;
        RECT 146.575 104.890 148.275 106.290 ;
        RECT 148.575 104.890 150.275 106.290 ;
        RECT 150.575 104.890 152.275 106.290 ;
        RECT 152.575 104.890 154.275 106.290 ;
        RECT 6.840 103.040 8.540 104.440 ;
        RECT 8.840 103.040 10.540 104.440 ;
        RECT 10.840 103.040 12.540 104.440 ;
        RECT 12.840 103.040 14.540 104.440 ;
        RECT 14.840 103.040 16.540 104.440 ;
        RECT 16.840 103.040 18.540 104.440 ;
        RECT 18.840 103.040 20.540 104.440 ;
        RECT 20.840 103.040 22.540 104.440 ;
        RECT 22.840 103.040 24.540 104.440 ;
        RECT 24.840 103.040 26.540 104.440 ;
        RECT 26.840 103.040 28.540 104.440 ;
        RECT 28.840 103.040 30.540 104.440 ;
        RECT 30.840 103.040 32.540 104.440 ;
        RECT 32.840 103.040 34.540 104.440 ;
        RECT 34.840 103.040 36.540 104.440 ;
        RECT 36.840 103.040 38.540 104.440 ;
        RECT 38.840 103.040 40.540 104.440 ;
        RECT 40.840 103.040 42.540 104.440 ;
        RECT 42.840 103.040 44.540 104.440 ;
        RECT 44.840 103.040 46.540 104.440 ;
        RECT 46.840 103.040 48.540 104.440 ;
        RECT 48.840 103.040 50.540 104.440 ;
        RECT 50.840 103.040 52.540 104.440 ;
        RECT 52.840 103.040 54.540 104.440 ;
        RECT 54.840 103.040 56.540 104.440 ;
        RECT 56.840 103.040 58.540 104.440 ;
        RECT 58.840 103.040 60.540 104.440 ;
        RECT 60.840 103.040 62.540 104.440 ;
        RECT 62.840 103.040 64.540 104.440 ;
        RECT 64.840 103.040 66.540 104.440 ;
        RECT 66.840 103.040 68.540 104.440 ;
        RECT 68.840 103.040 70.540 104.440 ;
        RECT 70.840 103.040 72.540 104.440 ;
        RECT 72.840 103.040 74.540 104.440 ;
        RECT 86.575 103.040 88.275 104.440 ;
        RECT 88.575 103.040 90.275 104.440 ;
        RECT 90.575 103.040 92.275 104.440 ;
        RECT 92.575 103.040 94.275 104.440 ;
        RECT 94.575 103.040 96.275 104.440 ;
        RECT 96.575 103.040 98.275 104.440 ;
        RECT 98.575 103.040 100.275 104.440 ;
        RECT 100.575 103.040 102.275 104.440 ;
        RECT 102.575 103.040 104.275 104.440 ;
        RECT 104.575 103.040 106.275 104.440 ;
        RECT 106.575 103.040 108.275 104.440 ;
        RECT 108.575 103.040 110.275 104.440 ;
        RECT 110.575 103.040 112.275 104.440 ;
        RECT 112.575 103.040 114.275 104.440 ;
        RECT 114.575 103.040 116.275 104.440 ;
        RECT 116.575 103.040 118.275 104.440 ;
        RECT 118.575 103.040 120.275 104.440 ;
        RECT 120.575 103.040 122.275 104.440 ;
        RECT 122.575 103.040 124.275 104.440 ;
        RECT 124.575 103.040 126.275 104.440 ;
        RECT 126.575 103.040 128.275 104.440 ;
        RECT 128.575 103.040 130.275 104.440 ;
        RECT 130.575 103.040 132.275 104.440 ;
        RECT 132.575 103.040 134.275 104.440 ;
        RECT 134.575 103.040 136.275 104.440 ;
        RECT 136.575 103.040 138.275 104.440 ;
        RECT 138.575 103.040 140.275 104.440 ;
        RECT 140.575 103.040 142.275 104.440 ;
        RECT 142.575 103.040 144.275 104.440 ;
        RECT 144.575 103.040 146.275 104.440 ;
        RECT 146.575 103.040 148.275 104.440 ;
        RECT 148.575 103.040 150.275 104.440 ;
        RECT 150.575 103.040 152.275 104.440 ;
        RECT 152.575 103.040 154.275 104.440 ;
        RECT 6.840 101.190 8.540 102.590 ;
        RECT 8.840 101.190 10.540 102.590 ;
        RECT 10.840 101.190 12.540 102.590 ;
        RECT 12.840 101.190 14.540 102.590 ;
        RECT 14.840 101.190 16.540 102.590 ;
        RECT 16.840 101.190 18.540 102.590 ;
        RECT 18.840 101.190 20.540 102.590 ;
        RECT 20.840 101.190 22.540 102.590 ;
        RECT 22.840 101.190 24.540 102.590 ;
        RECT 24.840 101.190 26.540 102.590 ;
        RECT 26.840 101.190 28.540 102.590 ;
        RECT 28.840 101.190 30.540 102.590 ;
        RECT 30.840 101.190 32.540 102.590 ;
        RECT 32.840 101.190 34.540 102.590 ;
        RECT 34.840 101.190 36.540 102.590 ;
        RECT 36.840 101.190 38.540 102.590 ;
        RECT 38.840 101.190 40.540 102.590 ;
        RECT 40.840 101.190 42.540 102.590 ;
        RECT 42.840 101.190 44.540 102.590 ;
        RECT 44.840 101.190 46.540 102.590 ;
        RECT 46.840 101.190 48.540 102.590 ;
        RECT 48.840 101.190 50.540 102.590 ;
        RECT 50.840 101.190 52.540 102.590 ;
        RECT 52.840 101.190 54.540 102.590 ;
        RECT 54.840 101.190 56.540 102.590 ;
        RECT 56.840 101.190 58.540 102.590 ;
        RECT 58.840 101.190 60.540 102.590 ;
        RECT 60.840 101.190 62.540 102.590 ;
        RECT 62.840 101.190 64.540 102.590 ;
        RECT 64.840 101.190 66.540 102.590 ;
        RECT 66.840 101.190 68.540 102.590 ;
        RECT 68.840 101.190 70.540 102.590 ;
        RECT 70.840 101.190 72.540 102.590 ;
        RECT 72.840 101.190 74.540 102.590 ;
        RECT 86.575 101.190 88.275 102.590 ;
        RECT 88.575 101.190 90.275 102.590 ;
        RECT 90.575 101.190 92.275 102.590 ;
        RECT 92.575 101.190 94.275 102.590 ;
        RECT 94.575 101.190 96.275 102.590 ;
        RECT 96.575 101.190 98.275 102.590 ;
        RECT 98.575 101.190 100.275 102.590 ;
        RECT 100.575 101.190 102.275 102.590 ;
        RECT 102.575 101.190 104.275 102.590 ;
        RECT 104.575 101.190 106.275 102.590 ;
        RECT 106.575 101.190 108.275 102.590 ;
        RECT 108.575 101.190 110.275 102.590 ;
        RECT 110.575 101.190 112.275 102.590 ;
        RECT 112.575 101.190 114.275 102.590 ;
        RECT 114.575 101.190 116.275 102.590 ;
        RECT 116.575 101.190 118.275 102.590 ;
        RECT 118.575 101.190 120.275 102.590 ;
        RECT 120.575 101.190 122.275 102.590 ;
        RECT 122.575 101.190 124.275 102.590 ;
        RECT 124.575 101.190 126.275 102.590 ;
        RECT 126.575 101.190 128.275 102.590 ;
        RECT 128.575 101.190 130.275 102.590 ;
        RECT 130.575 101.190 132.275 102.590 ;
        RECT 132.575 101.190 134.275 102.590 ;
        RECT 134.575 101.190 136.275 102.590 ;
        RECT 136.575 101.190 138.275 102.590 ;
        RECT 138.575 101.190 140.275 102.590 ;
        RECT 140.575 101.190 142.275 102.590 ;
        RECT 142.575 101.190 144.275 102.590 ;
        RECT 144.575 101.190 146.275 102.590 ;
        RECT 146.575 101.190 148.275 102.590 ;
        RECT 148.575 101.190 150.275 102.590 ;
        RECT 150.575 101.190 152.275 102.590 ;
        RECT 152.575 101.190 154.275 102.590 ;
        RECT 6.840 99.340 8.540 100.740 ;
        RECT 8.840 99.340 10.540 100.740 ;
        RECT 10.840 99.340 12.540 100.740 ;
        RECT 12.840 99.340 14.540 100.740 ;
        RECT 14.840 99.340 16.540 100.740 ;
        RECT 16.840 99.340 18.540 100.740 ;
        RECT 18.840 99.340 20.540 100.740 ;
        RECT 20.840 99.340 22.540 100.740 ;
        RECT 22.840 99.340 24.540 100.740 ;
        RECT 24.840 99.340 26.540 100.740 ;
        RECT 26.840 99.340 28.540 100.740 ;
        RECT 28.840 99.340 30.540 100.740 ;
        RECT 30.840 99.340 32.540 100.740 ;
        RECT 32.840 99.340 34.540 100.740 ;
        RECT 34.840 99.340 36.540 100.740 ;
        RECT 36.840 99.340 38.540 100.740 ;
        RECT 38.840 99.340 40.540 100.740 ;
        RECT 40.840 99.340 42.540 100.740 ;
        RECT 42.840 99.340 44.540 100.740 ;
        RECT 44.840 99.340 46.540 100.740 ;
        RECT 46.840 99.340 48.540 100.740 ;
        RECT 48.840 99.340 50.540 100.740 ;
        RECT 50.840 99.340 52.540 100.740 ;
        RECT 52.840 99.340 54.540 100.740 ;
        RECT 54.840 99.340 56.540 100.740 ;
        RECT 56.840 99.340 58.540 100.740 ;
        RECT 58.840 99.340 60.540 100.740 ;
        RECT 60.840 99.340 62.540 100.740 ;
        RECT 62.840 99.340 64.540 100.740 ;
        RECT 64.840 99.340 66.540 100.740 ;
        RECT 66.840 99.340 68.540 100.740 ;
        RECT 68.840 99.340 70.540 100.740 ;
        RECT 70.840 99.340 72.540 100.740 ;
        RECT 72.840 99.340 74.540 100.740 ;
        RECT 86.575 99.340 88.275 100.740 ;
        RECT 88.575 99.340 90.275 100.740 ;
        RECT 90.575 99.340 92.275 100.740 ;
        RECT 92.575 99.340 94.275 100.740 ;
        RECT 94.575 99.340 96.275 100.740 ;
        RECT 96.575 99.340 98.275 100.740 ;
        RECT 98.575 99.340 100.275 100.740 ;
        RECT 100.575 99.340 102.275 100.740 ;
        RECT 102.575 99.340 104.275 100.740 ;
        RECT 104.575 99.340 106.275 100.740 ;
        RECT 106.575 99.340 108.275 100.740 ;
        RECT 108.575 99.340 110.275 100.740 ;
        RECT 110.575 99.340 112.275 100.740 ;
        RECT 112.575 99.340 114.275 100.740 ;
        RECT 114.575 99.340 116.275 100.740 ;
        RECT 116.575 99.340 118.275 100.740 ;
        RECT 118.575 99.340 120.275 100.740 ;
        RECT 120.575 99.340 122.275 100.740 ;
        RECT 122.575 99.340 124.275 100.740 ;
        RECT 124.575 99.340 126.275 100.740 ;
        RECT 126.575 99.340 128.275 100.740 ;
        RECT 128.575 99.340 130.275 100.740 ;
        RECT 130.575 99.340 132.275 100.740 ;
        RECT 132.575 99.340 134.275 100.740 ;
        RECT 134.575 99.340 136.275 100.740 ;
        RECT 136.575 99.340 138.275 100.740 ;
        RECT 138.575 99.340 140.275 100.740 ;
        RECT 140.575 99.340 142.275 100.740 ;
        RECT 142.575 99.340 144.275 100.740 ;
        RECT 144.575 99.340 146.275 100.740 ;
        RECT 146.575 99.340 148.275 100.740 ;
        RECT 148.575 99.340 150.275 100.740 ;
        RECT 150.575 99.340 152.275 100.740 ;
        RECT 152.575 99.340 154.275 100.740 ;
        RECT 6.840 97.490 8.540 98.890 ;
        RECT 8.840 97.490 10.540 98.890 ;
        RECT 10.840 97.490 12.540 98.890 ;
        RECT 12.840 97.490 14.540 98.890 ;
        RECT 14.840 97.490 16.540 98.890 ;
        RECT 16.840 97.490 18.540 98.890 ;
        RECT 18.840 97.490 20.540 98.890 ;
        RECT 20.840 97.490 22.540 98.890 ;
        RECT 22.840 97.490 24.540 98.890 ;
        RECT 24.840 97.490 26.540 98.890 ;
        RECT 26.840 97.490 28.540 98.890 ;
        RECT 28.840 97.490 30.540 98.890 ;
        RECT 30.840 97.490 32.540 98.890 ;
        RECT 32.840 97.490 34.540 98.890 ;
        RECT 34.840 97.490 36.540 98.890 ;
        RECT 36.840 97.490 38.540 98.890 ;
        RECT 38.840 97.490 40.540 98.890 ;
        RECT 40.840 97.490 42.540 98.890 ;
        RECT 42.840 97.490 44.540 98.890 ;
        RECT 44.840 97.490 46.540 98.890 ;
        RECT 46.840 97.490 48.540 98.890 ;
        RECT 48.840 97.490 50.540 98.890 ;
        RECT 50.840 97.490 52.540 98.890 ;
        RECT 52.840 97.490 54.540 98.890 ;
        RECT 54.840 97.490 56.540 98.890 ;
        RECT 56.840 97.490 58.540 98.890 ;
        RECT 58.840 97.490 60.540 98.890 ;
        RECT 60.840 97.490 62.540 98.890 ;
        RECT 62.840 97.490 64.540 98.890 ;
        RECT 64.840 97.490 66.540 98.890 ;
        RECT 66.840 97.490 68.540 98.890 ;
        RECT 68.840 97.490 70.540 98.890 ;
        RECT 70.840 97.490 72.540 98.890 ;
        RECT 72.840 97.490 74.540 98.890 ;
        RECT 86.575 97.490 88.275 98.890 ;
        RECT 88.575 97.490 90.275 98.890 ;
        RECT 90.575 97.490 92.275 98.890 ;
        RECT 92.575 97.490 94.275 98.890 ;
        RECT 94.575 97.490 96.275 98.890 ;
        RECT 96.575 97.490 98.275 98.890 ;
        RECT 98.575 97.490 100.275 98.890 ;
        RECT 100.575 97.490 102.275 98.890 ;
        RECT 102.575 97.490 104.275 98.890 ;
        RECT 104.575 97.490 106.275 98.890 ;
        RECT 106.575 97.490 108.275 98.890 ;
        RECT 108.575 97.490 110.275 98.890 ;
        RECT 110.575 97.490 112.275 98.890 ;
        RECT 112.575 97.490 114.275 98.890 ;
        RECT 114.575 97.490 116.275 98.890 ;
        RECT 116.575 97.490 118.275 98.890 ;
        RECT 118.575 97.490 120.275 98.890 ;
        RECT 120.575 97.490 122.275 98.890 ;
        RECT 122.575 97.490 124.275 98.890 ;
        RECT 124.575 97.490 126.275 98.890 ;
        RECT 126.575 97.490 128.275 98.890 ;
        RECT 128.575 97.490 130.275 98.890 ;
        RECT 130.575 97.490 132.275 98.890 ;
        RECT 132.575 97.490 134.275 98.890 ;
        RECT 134.575 97.490 136.275 98.890 ;
        RECT 136.575 97.490 138.275 98.890 ;
        RECT 138.575 97.490 140.275 98.890 ;
        RECT 140.575 97.490 142.275 98.890 ;
        RECT 142.575 97.490 144.275 98.890 ;
        RECT 144.575 97.490 146.275 98.890 ;
        RECT 146.575 97.490 148.275 98.890 ;
        RECT 148.575 97.490 150.275 98.890 ;
        RECT 150.575 97.490 152.275 98.890 ;
        RECT 152.575 97.490 154.275 98.890 ;
        RECT 6.840 95.640 8.540 97.040 ;
        RECT 8.840 95.640 10.540 97.040 ;
        RECT 10.840 95.640 12.540 97.040 ;
        RECT 12.840 95.640 14.540 97.040 ;
        RECT 14.840 95.640 16.540 97.040 ;
        RECT 16.840 95.640 18.540 97.040 ;
        RECT 18.840 95.640 20.540 97.040 ;
        RECT 20.840 95.640 22.540 97.040 ;
        RECT 22.840 95.640 24.540 97.040 ;
        RECT 24.840 95.640 26.540 97.040 ;
        RECT 26.840 95.640 28.540 97.040 ;
        RECT 28.840 95.640 30.540 97.040 ;
        RECT 30.840 95.640 32.540 97.040 ;
        RECT 32.840 95.640 34.540 97.040 ;
        RECT 34.840 95.640 36.540 97.040 ;
        RECT 36.840 95.640 38.540 97.040 ;
        RECT 38.840 95.640 40.540 97.040 ;
        RECT 40.840 95.640 42.540 97.040 ;
        RECT 42.840 95.640 44.540 97.040 ;
        RECT 44.840 95.640 46.540 97.040 ;
        RECT 46.840 95.640 48.540 97.040 ;
        RECT 48.840 95.640 50.540 97.040 ;
        RECT 50.840 95.640 52.540 97.040 ;
        RECT 52.840 95.640 54.540 97.040 ;
        RECT 54.840 95.640 56.540 97.040 ;
        RECT 56.840 95.640 58.540 97.040 ;
        RECT 58.840 95.640 60.540 97.040 ;
        RECT 60.840 95.640 62.540 97.040 ;
        RECT 62.840 95.640 64.540 97.040 ;
        RECT 64.840 95.640 66.540 97.040 ;
        RECT 66.840 95.640 68.540 97.040 ;
        RECT 68.840 95.640 70.540 97.040 ;
        RECT 70.840 95.640 72.540 97.040 ;
        RECT 72.840 95.640 74.540 97.040 ;
        RECT 86.575 95.640 88.275 97.040 ;
        RECT 88.575 95.640 90.275 97.040 ;
        RECT 90.575 95.640 92.275 97.040 ;
        RECT 92.575 95.640 94.275 97.040 ;
        RECT 94.575 95.640 96.275 97.040 ;
        RECT 96.575 95.640 98.275 97.040 ;
        RECT 98.575 95.640 100.275 97.040 ;
        RECT 100.575 95.640 102.275 97.040 ;
        RECT 102.575 95.640 104.275 97.040 ;
        RECT 104.575 95.640 106.275 97.040 ;
        RECT 106.575 95.640 108.275 97.040 ;
        RECT 108.575 95.640 110.275 97.040 ;
        RECT 110.575 95.640 112.275 97.040 ;
        RECT 112.575 95.640 114.275 97.040 ;
        RECT 114.575 95.640 116.275 97.040 ;
        RECT 116.575 95.640 118.275 97.040 ;
        RECT 118.575 95.640 120.275 97.040 ;
        RECT 120.575 95.640 122.275 97.040 ;
        RECT 122.575 95.640 124.275 97.040 ;
        RECT 124.575 95.640 126.275 97.040 ;
        RECT 126.575 95.640 128.275 97.040 ;
        RECT 128.575 95.640 130.275 97.040 ;
        RECT 130.575 95.640 132.275 97.040 ;
        RECT 132.575 95.640 134.275 97.040 ;
        RECT 134.575 95.640 136.275 97.040 ;
        RECT 136.575 95.640 138.275 97.040 ;
        RECT 138.575 95.640 140.275 97.040 ;
        RECT 140.575 95.640 142.275 97.040 ;
        RECT 142.575 95.640 144.275 97.040 ;
        RECT 144.575 95.640 146.275 97.040 ;
        RECT 146.575 95.640 148.275 97.040 ;
        RECT 148.575 95.640 150.275 97.040 ;
        RECT 150.575 95.640 152.275 97.040 ;
        RECT 152.575 95.640 154.275 97.040 ;
        RECT 6.840 93.790 8.540 95.190 ;
        RECT 8.840 93.790 10.540 95.190 ;
        RECT 10.840 93.790 12.540 95.190 ;
        RECT 12.840 93.790 14.540 95.190 ;
        RECT 14.840 93.790 16.540 95.190 ;
        RECT 16.840 93.790 18.540 95.190 ;
        RECT 18.840 93.790 20.540 95.190 ;
        RECT 20.840 93.790 22.540 95.190 ;
        RECT 22.840 93.790 24.540 95.190 ;
        RECT 24.840 93.790 26.540 95.190 ;
        RECT 26.840 93.790 28.540 95.190 ;
        RECT 28.840 93.790 30.540 95.190 ;
        RECT 30.840 93.790 32.540 95.190 ;
        RECT 32.840 93.790 34.540 95.190 ;
        RECT 34.840 93.790 36.540 95.190 ;
        RECT 36.840 93.790 38.540 95.190 ;
        RECT 38.840 93.790 40.540 95.190 ;
        RECT 40.840 93.790 42.540 95.190 ;
        RECT 42.840 93.790 44.540 95.190 ;
        RECT 44.840 93.790 46.540 95.190 ;
        RECT 46.840 93.790 48.540 95.190 ;
        RECT 48.840 93.790 50.540 95.190 ;
        RECT 50.840 93.790 52.540 95.190 ;
        RECT 52.840 93.790 54.540 95.190 ;
        RECT 54.840 93.790 56.540 95.190 ;
        RECT 56.840 93.790 58.540 95.190 ;
        RECT 58.840 93.790 60.540 95.190 ;
        RECT 60.840 93.790 62.540 95.190 ;
        RECT 62.840 93.790 64.540 95.190 ;
        RECT 64.840 93.790 66.540 95.190 ;
        RECT 66.840 93.790 68.540 95.190 ;
        RECT 68.840 93.790 70.540 95.190 ;
        RECT 70.840 93.790 72.540 95.190 ;
        RECT 72.840 93.790 74.540 95.190 ;
        RECT 86.575 93.790 88.275 95.190 ;
        RECT 88.575 93.790 90.275 95.190 ;
        RECT 90.575 93.790 92.275 95.190 ;
        RECT 92.575 93.790 94.275 95.190 ;
        RECT 94.575 93.790 96.275 95.190 ;
        RECT 96.575 93.790 98.275 95.190 ;
        RECT 98.575 93.790 100.275 95.190 ;
        RECT 100.575 93.790 102.275 95.190 ;
        RECT 102.575 93.790 104.275 95.190 ;
        RECT 104.575 93.790 106.275 95.190 ;
        RECT 106.575 93.790 108.275 95.190 ;
        RECT 108.575 93.790 110.275 95.190 ;
        RECT 110.575 93.790 112.275 95.190 ;
        RECT 112.575 93.790 114.275 95.190 ;
        RECT 114.575 93.790 116.275 95.190 ;
        RECT 116.575 93.790 118.275 95.190 ;
        RECT 118.575 93.790 120.275 95.190 ;
        RECT 120.575 93.790 122.275 95.190 ;
        RECT 122.575 93.790 124.275 95.190 ;
        RECT 124.575 93.790 126.275 95.190 ;
        RECT 126.575 93.790 128.275 95.190 ;
        RECT 128.575 93.790 130.275 95.190 ;
        RECT 130.575 93.790 132.275 95.190 ;
        RECT 132.575 93.790 134.275 95.190 ;
        RECT 134.575 93.790 136.275 95.190 ;
        RECT 136.575 93.790 138.275 95.190 ;
        RECT 138.575 93.790 140.275 95.190 ;
        RECT 140.575 93.790 142.275 95.190 ;
        RECT 142.575 93.790 144.275 95.190 ;
        RECT 144.575 93.790 146.275 95.190 ;
        RECT 146.575 93.790 148.275 95.190 ;
        RECT 148.575 93.790 150.275 95.190 ;
        RECT 150.575 93.790 152.275 95.190 ;
        RECT 152.575 93.790 154.275 95.190 ;
        RECT 6.840 91.940 8.540 93.340 ;
        RECT 8.840 91.940 10.540 93.340 ;
        RECT 10.840 91.940 12.540 93.340 ;
        RECT 12.840 91.940 14.540 93.340 ;
        RECT 14.840 91.940 16.540 93.340 ;
        RECT 16.840 91.940 18.540 93.340 ;
        RECT 18.840 91.940 20.540 93.340 ;
        RECT 20.840 91.940 22.540 93.340 ;
        RECT 22.840 91.940 24.540 93.340 ;
        RECT 24.840 91.940 26.540 93.340 ;
        RECT 26.840 91.940 28.540 93.340 ;
        RECT 28.840 91.940 30.540 93.340 ;
        RECT 30.840 91.940 32.540 93.340 ;
        RECT 32.840 91.940 34.540 93.340 ;
        RECT 34.840 91.940 36.540 93.340 ;
        RECT 36.840 91.940 38.540 93.340 ;
        RECT 38.840 91.940 40.540 93.340 ;
        RECT 40.840 91.940 42.540 93.340 ;
        RECT 42.840 91.940 44.540 93.340 ;
        RECT 44.840 91.940 46.540 93.340 ;
        RECT 46.840 91.940 48.540 93.340 ;
        RECT 48.840 91.940 50.540 93.340 ;
        RECT 50.840 91.940 52.540 93.340 ;
        RECT 52.840 91.940 54.540 93.340 ;
        RECT 54.840 91.940 56.540 93.340 ;
        RECT 56.840 91.940 58.540 93.340 ;
        RECT 58.840 91.940 60.540 93.340 ;
        RECT 60.840 91.940 62.540 93.340 ;
        RECT 62.840 91.940 64.540 93.340 ;
        RECT 64.840 91.940 66.540 93.340 ;
        RECT 66.840 91.940 68.540 93.340 ;
        RECT 68.840 91.940 70.540 93.340 ;
        RECT 70.840 91.940 72.540 93.340 ;
        RECT 72.840 91.940 74.540 93.340 ;
        RECT 86.575 91.940 88.275 93.340 ;
        RECT 88.575 91.940 90.275 93.340 ;
        RECT 90.575 91.940 92.275 93.340 ;
        RECT 92.575 91.940 94.275 93.340 ;
        RECT 94.575 91.940 96.275 93.340 ;
        RECT 96.575 91.940 98.275 93.340 ;
        RECT 98.575 91.940 100.275 93.340 ;
        RECT 100.575 91.940 102.275 93.340 ;
        RECT 102.575 91.940 104.275 93.340 ;
        RECT 104.575 91.940 106.275 93.340 ;
        RECT 106.575 91.940 108.275 93.340 ;
        RECT 108.575 91.940 110.275 93.340 ;
        RECT 110.575 91.940 112.275 93.340 ;
        RECT 112.575 91.940 114.275 93.340 ;
        RECT 114.575 91.940 116.275 93.340 ;
        RECT 116.575 91.940 118.275 93.340 ;
        RECT 118.575 91.940 120.275 93.340 ;
        RECT 120.575 91.940 122.275 93.340 ;
        RECT 122.575 91.940 124.275 93.340 ;
        RECT 124.575 91.940 126.275 93.340 ;
        RECT 126.575 91.940 128.275 93.340 ;
        RECT 128.575 91.940 130.275 93.340 ;
        RECT 130.575 91.940 132.275 93.340 ;
        RECT 132.575 91.940 134.275 93.340 ;
        RECT 134.575 91.940 136.275 93.340 ;
        RECT 136.575 91.940 138.275 93.340 ;
        RECT 138.575 91.940 140.275 93.340 ;
        RECT 140.575 91.940 142.275 93.340 ;
        RECT 142.575 91.940 144.275 93.340 ;
        RECT 144.575 91.940 146.275 93.340 ;
        RECT 146.575 91.940 148.275 93.340 ;
        RECT 148.575 91.940 150.275 93.340 ;
        RECT 150.575 91.940 152.275 93.340 ;
        RECT 152.575 91.940 154.275 93.340 ;
        RECT 6.840 90.090 8.540 91.490 ;
        RECT 8.840 90.090 10.540 91.490 ;
        RECT 10.840 90.090 12.540 91.490 ;
        RECT 12.840 90.090 14.540 91.490 ;
        RECT 14.840 90.090 16.540 91.490 ;
        RECT 16.840 90.090 18.540 91.490 ;
        RECT 18.840 90.090 20.540 91.490 ;
        RECT 20.840 90.090 22.540 91.490 ;
        RECT 22.840 90.090 24.540 91.490 ;
        RECT 24.840 90.090 26.540 91.490 ;
        RECT 26.840 90.090 28.540 91.490 ;
        RECT 28.840 90.090 30.540 91.490 ;
        RECT 30.840 90.090 32.540 91.490 ;
        RECT 32.840 90.090 34.540 91.490 ;
        RECT 34.840 90.090 36.540 91.490 ;
        RECT 36.840 90.090 38.540 91.490 ;
        RECT 38.840 90.090 40.540 91.490 ;
        RECT 40.840 90.090 42.540 91.490 ;
        RECT 42.840 90.090 44.540 91.490 ;
        RECT 44.840 90.090 46.540 91.490 ;
        RECT 46.840 90.090 48.540 91.490 ;
        RECT 48.840 90.090 50.540 91.490 ;
        RECT 50.840 90.090 52.540 91.490 ;
        RECT 52.840 90.090 54.540 91.490 ;
        RECT 54.840 90.090 56.540 91.490 ;
        RECT 56.840 90.090 58.540 91.490 ;
        RECT 58.840 90.090 60.540 91.490 ;
        RECT 60.840 90.090 62.540 91.490 ;
        RECT 62.840 90.090 64.540 91.490 ;
        RECT 64.840 90.090 66.540 91.490 ;
        RECT 66.840 90.090 68.540 91.490 ;
        RECT 68.840 90.090 70.540 91.490 ;
        RECT 70.840 90.090 72.540 91.490 ;
        RECT 72.840 90.090 74.540 91.490 ;
        RECT 86.575 90.090 88.275 91.490 ;
        RECT 88.575 90.090 90.275 91.490 ;
        RECT 90.575 90.090 92.275 91.490 ;
        RECT 92.575 90.090 94.275 91.490 ;
        RECT 94.575 90.090 96.275 91.490 ;
        RECT 96.575 90.090 98.275 91.490 ;
        RECT 98.575 90.090 100.275 91.490 ;
        RECT 100.575 90.090 102.275 91.490 ;
        RECT 102.575 90.090 104.275 91.490 ;
        RECT 104.575 90.090 106.275 91.490 ;
        RECT 106.575 90.090 108.275 91.490 ;
        RECT 108.575 90.090 110.275 91.490 ;
        RECT 110.575 90.090 112.275 91.490 ;
        RECT 112.575 90.090 114.275 91.490 ;
        RECT 114.575 90.090 116.275 91.490 ;
        RECT 116.575 90.090 118.275 91.490 ;
        RECT 118.575 90.090 120.275 91.490 ;
        RECT 120.575 90.090 122.275 91.490 ;
        RECT 122.575 90.090 124.275 91.490 ;
        RECT 124.575 90.090 126.275 91.490 ;
        RECT 126.575 90.090 128.275 91.490 ;
        RECT 128.575 90.090 130.275 91.490 ;
        RECT 130.575 90.090 132.275 91.490 ;
        RECT 132.575 90.090 134.275 91.490 ;
        RECT 134.575 90.090 136.275 91.490 ;
        RECT 136.575 90.090 138.275 91.490 ;
        RECT 138.575 90.090 140.275 91.490 ;
        RECT 140.575 90.090 142.275 91.490 ;
        RECT 142.575 90.090 144.275 91.490 ;
        RECT 144.575 90.090 146.275 91.490 ;
        RECT 146.575 90.090 148.275 91.490 ;
        RECT 148.575 90.090 150.275 91.490 ;
        RECT 150.575 90.090 152.275 91.490 ;
        RECT 152.575 90.090 154.275 91.490 ;
        RECT 6.840 88.240 8.540 89.640 ;
        RECT 8.840 88.240 10.540 89.640 ;
        RECT 10.840 88.240 12.540 89.640 ;
        RECT 12.840 88.240 14.540 89.640 ;
        RECT 14.840 88.240 16.540 89.640 ;
        RECT 16.840 88.240 18.540 89.640 ;
        RECT 18.840 88.240 20.540 89.640 ;
        RECT 20.840 88.240 22.540 89.640 ;
        RECT 22.840 88.240 24.540 89.640 ;
        RECT 24.840 88.240 26.540 89.640 ;
        RECT 26.840 88.240 28.540 89.640 ;
        RECT 28.840 88.240 30.540 89.640 ;
        RECT 30.840 88.240 32.540 89.640 ;
        RECT 32.840 88.240 34.540 89.640 ;
        RECT 34.840 88.240 36.540 89.640 ;
        RECT 36.840 88.240 38.540 89.640 ;
        RECT 38.840 88.240 40.540 89.640 ;
        RECT 40.840 88.240 42.540 89.640 ;
        RECT 42.840 88.240 44.540 89.640 ;
        RECT 44.840 88.240 46.540 89.640 ;
        RECT 46.840 88.240 48.540 89.640 ;
        RECT 48.840 88.240 50.540 89.640 ;
        RECT 50.840 88.240 52.540 89.640 ;
        RECT 52.840 88.240 54.540 89.640 ;
        RECT 54.840 88.240 56.540 89.640 ;
        RECT 56.840 88.240 58.540 89.640 ;
        RECT 58.840 88.240 60.540 89.640 ;
        RECT 60.840 88.240 62.540 89.640 ;
        RECT 62.840 88.240 64.540 89.640 ;
        RECT 64.840 88.240 66.540 89.640 ;
        RECT 66.840 88.240 68.540 89.640 ;
        RECT 68.840 88.240 70.540 89.640 ;
        RECT 70.840 88.240 72.540 89.640 ;
        RECT 72.840 88.240 74.540 89.640 ;
        RECT 86.575 88.240 88.275 89.640 ;
        RECT 88.575 88.240 90.275 89.640 ;
        RECT 90.575 88.240 92.275 89.640 ;
        RECT 92.575 88.240 94.275 89.640 ;
        RECT 94.575 88.240 96.275 89.640 ;
        RECT 96.575 88.240 98.275 89.640 ;
        RECT 98.575 88.240 100.275 89.640 ;
        RECT 100.575 88.240 102.275 89.640 ;
        RECT 102.575 88.240 104.275 89.640 ;
        RECT 104.575 88.240 106.275 89.640 ;
        RECT 106.575 88.240 108.275 89.640 ;
        RECT 108.575 88.240 110.275 89.640 ;
        RECT 110.575 88.240 112.275 89.640 ;
        RECT 112.575 88.240 114.275 89.640 ;
        RECT 114.575 88.240 116.275 89.640 ;
        RECT 116.575 88.240 118.275 89.640 ;
        RECT 118.575 88.240 120.275 89.640 ;
        RECT 120.575 88.240 122.275 89.640 ;
        RECT 122.575 88.240 124.275 89.640 ;
        RECT 124.575 88.240 126.275 89.640 ;
        RECT 126.575 88.240 128.275 89.640 ;
        RECT 128.575 88.240 130.275 89.640 ;
        RECT 130.575 88.240 132.275 89.640 ;
        RECT 132.575 88.240 134.275 89.640 ;
        RECT 134.575 88.240 136.275 89.640 ;
        RECT 136.575 88.240 138.275 89.640 ;
        RECT 138.575 88.240 140.275 89.640 ;
        RECT 140.575 88.240 142.275 89.640 ;
        RECT 142.575 88.240 144.275 89.640 ;
        RECT 144.575 88.240 146.275 89.640 ;
        RECT 146.575 88.240 148.275 89.640 ;
        RECT 148.575 88.240 150.275 89.640 ;
        RECT 150.575 88.240 152.275 89.640 ;
        RECT 152.575 88.240 154.275 89.640 ;
        RECT 6.840 86.390 8.540 87.790 ;
        RECT 8.840 86.390 10.540 87.790 ;
        RECT 10.840 86.390 12.540 87.790 ;
        RECT 12.840 86.390 14.540 87.790 ;
        RECT 14.840 86.390 16.540 87.790 ;
        RECT 16.840 86.390 18.540 87.790 ;
        RECT 18.840 86.390 20.540 87.790 ;
        RECT 20.840 86.390 22.540 87.790 ;
        RECT 22.840 86.390 24.540 87.790 ;
        RECT 24.840 86.390 26.540 87.790 ;
        RECT 26.840 86.390 28.540 87.790 ;
        RECT 28.840 86.390 30.540 87.790 ;
        RECT 30.840 86.390 32.540 87.790 ;
        RECT 32.840 86.390 34.540 87.790 ;
        RECT 34.840 86.390 36.540 87.790 ;
        RECT 36.840 86.390 38.540 87.790 ;
        RECT 38.840 86.390 40.540 87.790 ;
        RECT 40.840 86.390 42.540 87.790 ;
        RECT 42.840 86.390 44.540 87.790 ;
        RECT 44.840 86.390 46.540 87.790 ;
        RECT 46.840 86.390 48.540 87.790 ;
        RECT 48.840 86.390 50.540 87.790 ;
        RECT 50.840 86.390 52.540 87.790 ;
        RECT 52.840 86.390 54.540 87.790 ;
        RECT 54.840 86.390 56.540 87.790 ;
        RECT 56.840 86.390 58.540 87.790 ;
        RECT 58.840 86.390 60.540 87.790 ;
        RECT 60.840 86.390 62.540 87.790 ;
        RECT 62.840 86.390 64.540 87.790 ;
        RECT 64.840 86.390 66.540 87.790 ;
        RECT 66.840 86.390 68.540 87.790 ;
        RECT 68.840 86.390 70.540 87.790 ;
        RECT 70.840 86.390 72.540 87.790 ;
        RECT 72.840 86.390 74.540 87.790 ;
        RECT 86.575 86.390 88.275 87.790 ;
        RECT 88.575 86.390 90.275 87.790 ;
        RECT 90.575 86.390 92.275 87.790 ;
        RECT 92.575 86.390 94.275 87.790 ;
        RECT 94.575 86.390 96.275 87.790 ;
        RECT 96.575 86.390 98.275 87.790 ;
        RECT 98.575 86.390 100.275 87.790 ;
        RECT 100.575 86.390 102.275 87.790 ;
        RECT 102.575 86.390 104.275 87.790 ;
        RECT 104.575 86.390 106.275 87.790 ;
        RECT 106.575 86.390 108.275 87.790 ;
        RECT 108.575 86.390 110.275 87.790 ;
        RECT 110.575 86.390 112.275 87.790 ;
        RECT 112.575 86.390 114.275 87.790 ;
        RECT 114.575 86.390 116.275 87.790 ;
        RECT 116.575 86.390 118.275 87.790 ;
        RECT 118.575 86.390 120.275 87.790 ;
        RECT 120.575 86.390 122.275 87.790 ;
        RECT 122.575 86.390 124.275 87.790 ;
        RECT 124.575 86.390 126.275 87.790 ;
        RECT 126.575 86.390 128.275 87.790 ;
        RECT 128.575 86.390 130.275 87.790 ;
        RECT 130.575 86.390 132.275 87.790 ;
        RECT 132.575 86.390 134.275 87.790 ;
        RECT 134.575 86.390 136.275 87.790 ;
        RECT 136.575 86.390 138.275 87.790 ;
        RECT 138.575 86.390 140.275 87.790 ;
        RECT 140.575 86.390 142.275 87.790 ;
        RECT 142.575 86.390 144.275 87.790 ;
        RECT 144.575 86.390 146.275 87.790 ;
        RECT 146.575 86.390 148.275 87.790 ;
        RECT 148.575 86.390 150.275 87.790 ;
        RECT 150.575 86.390 152.275 87.790 ;
        RECT 152.575 86.390 154.275 87.790 ;
        RECT 6.840 84.540 8.540 85.940 ;
        RECT 8.840 84.540 10.540 85.940 ;
        RECT 10.840 84.540 12.540 85.940 ;
        RECT 12.840 84.540 14.540 85.940 ;
        RECT 14.840 84.540 16.540 85.940 ;
        RECT 16.840 84.540 18.540 85.940 ;
        RECT 18.840 84.540 20.540 85.940 ;
        RECT 20.840 84.540 22.540 85.940 ;
        RECT 22.840 84.540 24.540 85.940 ;
        RECT 24.840 84.540 26.540 85.940 ;
        RECT 26.840 84.540 28.540 85.940 ;
        RECT 28.840 84.540 30.540 85.940 ;
        RECT 30.840 84.540 32.540 85.940 ;
        RECT 32.840 84.540 34.540 85.940 ;
        RECT 34.840 84.540 36.540 85.940 ;
        RECT 36.840 84.540 38.540 85.940 ;
        RECT 38.840 84.540 40.540 85.940 ;
        RECT 40.840 84.540 42.540 85.940 ;
        RECT 42.840 84.540 44.540 85.940 ;
        RECT 44.840 84.540 46.540 85.940 ;
        RECT 46.840 84.540 48.540 85.940 ;
        RECT 48.840 84.540 50.540 85.940 ;
        RECT 50.840 84.540 52.540 85.940 ;
        RECT 52.840 84.540 54.540 85.940 ;
        RECT 54.840 84.540 56.540 85.940 ;
        RECT 56.840 84.540 58.540 85.940 ;
        RECT 58.840 84.540 60.540 85.940 ;
        RECT 60.840 84.540 62.540 85.940 ;
        RECT 62.840 84.540 64.540 85.940 ;
        RECT 64.840 84.540 66.540 85.940 ;
        RECT 66.840 84.540 68.540 85.940 ;
        RECT 68.840 84.540 70.540 85.940 ;
        RECT 70.840 84.540 72.540 85.940 ;
        RECT 72.840 84.540 74.540 85.940 ;
        RECT 86.575 84.540 88.275 85.940 ;
        RECT 88.575 84.540 90.275 85.940 ;
        RECT 90.575 84.540 92.275 85.940 ;
        RECT 92.575 84.540 94.275 85.940 ;
        RECT 94.575 84.540 96.275 85.940 ;
        RECT 96.575 84.540 98.275 85.940 ;
        RECT 98.575 84.540 100.275 85.940 ;
        RECT 100.575 84.540 102.275 85.940 ;
        RECT 102.575 84.540 104.275 85.940 ;
        RECT 104.575 84.540 106.275 85.940 ;
        RECT 106.575 84.540 108.275 85.940 ;
        RECT 108.575 84.540 110.275 85.940 ;
        RECT 110.575 84.540 112.275 85.940 ;
        RECT 112.575 84.540 114.275 85.940 ;
        RECT 114.575 84.540 116.275 85.940 ;
        RECT 116.575 84.540 118.275 85.940 ;
        RECT 118.575 84.540 120.275 85.940 ;
        RECT 120.575 84.540 122.275 85.940 ;
        RECT 122.575 84.540 124.275 85.940 ;
        RECT 124.575 84.540 126.275 85.940 ;
        RECT 126.575 84.540 128.275 85.940 ;
        RECT 128.575 84.540 130.275 85.940 ;
        RECT 130.575 84.540 132.275 85.940 ;
        RECT 132.575 84.540 134.275 85.940 ;
        RECT 134.575 84.540 136.275 85.940 ;
        RECT 136.575 84.540 138.275 85.940 ;
        RECT 138.575 84.540 140.275 85.940 ;
        RECT 140.575 84.540 142.275 85.940 ;
        RECT 142.575 84.540 144.275 85.940 ;
        RECT 144.575 84.540 146.275 85.940 ;
        RECT 146.575 84.540 148.275 85.940 ;
        RECT 148.575 84.540 150.275 85.940 ;
        RECT 150.575 84.540 152.275 85.940 ;
        RECT 152.575 84.540 154.275 85.940 ;
        RECT 6.840 82.690 8.540 84.090 ;
        RECT 8.840 82.690 10.540 84.090 ;
        RECT 10.840 82.690 12.540 84.090 ;
        RECT 12.840 82.690 14.540 84.090 ;
        RECT 14.840 82.690 16.540 84.090 ;
        RECT 16.840 82.690 18.540 84.090 ;
        RECT 18.840 82.690 20.540 84.090 ;
        RECT 20.840 82.690 22.540 84.090 ;
        RECT 22.840 82.690 24.540 84.090 ;
        RECT 24.840 82.690 26.540 84.090 ;
        RECT 26.840 82.690 28.540 84.090 ;
        RECT 28.840 82.690 30.540 84.090 ;
        RECT 30.840 82.690 32.540 84.090 ;
        RECT 32.840 82.690 34.540 84.090 ;
        RECT 34.840 82.690 36.540 84.090 ;
        RECT 36.840 82.690 38.540 84.090 ;
        RECT 38.840 82.690 40.540 84.090 ;
        RECT 40.840 82.690 42.540 84.090 ;
        RECT 42.840 82.690 44.540 84.090 ;
        RECT 44.840 82.690 46.540 84.090 ;
        RECT 46.840 82.690 48.540 84.090 ;
        RECT 48.840 82.690 50.540 84.090 ;
        RECT 50.840 82.690 52.540 84.090 ;
        RECT 52.840 82.690 54.540 84.090 ;
        RECT 54.840 82.690 56.540 84.090 ;
        RECT 56.840 82.690 58.540 84.090 ;
        RECT 58.840 82.690 60.540 84.090 ;
        RECT 60.840 82.690 62.540 84.090 ;
        RECT 62.840 82.690 64.540 84.090 ;
        RECT 64.840 82.690 66.540 84.090 ;
        RECT 66.840 82.690 68.540 84.090 ;
        RECT 68.840 82.690 70.540 84.090 ;
        RECT 70.840 82.690 72.540 84.090 ;
        RECT 72.840 82.690 74.540 84.090 ;
        RECT 86.575 82.690 88.275 84.090 ;
        RECT 88.575 82.690 90.275 84.090 ;
        RECT 90.575 82.690 92.275 84.090 ;
        RECT 92.575 82.690 94.275 84.090 ;
        RECT 94.575 82.690 96.275 84.090 ;
        RECT 96.575 82.690 98.275 84.090 ;
        RECT 98.575 82.690 100.275 84.090 ;
        RECT 100.575 82.690 102.275 84.090 ;
        RECT 102.575 82.690 104.275 84.090 ;
        RECT 104.575 82.690 106.275 84.090 ;
        RECT 106.575 82.690 108.275 84.090 ;
        RECT 108.575 82.690 110.275 84.090 ;
        RECT 110.575 82.690 112.275 84.090 ;
        RECT 112.575 82.690 114.275 84.090 ;
        RECT 114.575 82.690 116.275 84.090 ;
        RECT 116.575 82.690 118.275 84.090 ;
        RECT 118.575 82.690 120.275 84.090 ;
        RECT 120.575 82.690 122.275 84.090 ;
        RECT 122.575 82.690 124.275 84.090 ;
        RECT 124.575 82.690 126.275 84.090 ;
        RECT 126.575 82.690 128.275 84.090 ;
        RECT 128.575 82.690 130.275 84.090 ;
        RECT 130.575 82.690 132.275 84.090 ;
        RECT 132.575 82.690 134.275 84.090 ;
        RECT 134.575 82.690 136.275 84.090 ;
        RECT 136.575 82.690 138.275 84.090 ;
        RECT 138.575 82.690 140.275 84.090 ;
        RECT 140.575 82.690 142.275 84.090 ;
        RECT 142.575 82.690 144.275 84.090 ;
        RECT 144.575 82.690 146.275 84.090 ;
        RECT 146.575 82.690 148.275 84.090 ;
        RECT 148.575 82.690 150.275 84.090 ;
        RECT 150.575 82.690 152.275 84.090 ;
        RECT 152.575 82.690 154.275 84.090 ;
        RECT 6.840 80.840 8.540 82.240 ;
        RECT 8.840 80.840 10.540 82.240 ;
        RECT 10.840 80.840 12.540 82.240 ;
        RECT 12.840 80.840 14.540 82.240 ;
        RECT 14.840 80.840 16.540 82.240 ;
        RECT 16.840 80.840 18.540 82.240 ;
        RECT 18.840 80.840 20.540 82.240 ;
        RECT 20.840 80.840 22.540 82.240 ;
        RECT 22.840 80.840 24.540 82.240 ;
        RECT 24.840 80.840 26.540 82.240 ;
        RECT 26.840 80.840 28.540 82.240 ;
        RECT 28.840 80.840 30.540 82.240 ;
        RECT 30.840 80.840 32.540 82.240 ;
        RECT 32.840 80.840 34.540 82.240 ;
        RECT 34.840 80.840 36.540 82.240 ;
        RECT 36.840 80.840 38.540 82.240 ;
        RECT 38.840 80.840 40.540 82.240 ;
        RECT 40.840 80.840 42.540 82.240 ;
        RECT 42.840 80.840 44.540 82.240 ;
        RECT 44.840 80.840 46.540 82.240 ;
        RECT 46.840 80.840 48.540 82.240 ;
        RECT 48.840 80.840 50.540 82.240 ;
        RECT 50.840 80.840 52.540 82.240 ;
        RECT 52.840 80.840 54.540 82.240 ;
        RECT 54.840 80.840 56.540 82.240 ;
        RECT 56.840 80.840 58.540 82.240 ;
        RECT 58.840 80.840 60.540 82.240 ;
        RECT 60.840 80.840 62.540 82.240 ;
        RECT 62.840 80.840 64.540 82.240 ;
        RECT 64.840 80.840 66.540 82.240 ;
        RECT 66.840 80.840 68.540 82.240 ;
        RECT 68.840 80.840 70.540 82.240 ;
        RECT 70.840 80.840 72.540 82.240 ;
        RECT 72.840 80.840 74.540 82.240 ;
        RECT 86.575 80.840 88.275 82.240 ;
        RECT 88.575 80.840 90.275 82.240 ;
        RECT 90.575 80.840 92.275 82.240 ;
        RECT 92.575 80.840 94.275 82.240 ;
        RECT 94.575 80.840 96.275 82.240 ;
        RECT 96.575 80.840 98.275 82.240 ;
        RECT 98.575 80.840 100.275 82.240 ;
        RECT 100.575 80.840 102.275 82.240 ;
        RECT 102.575 80.840 104.275 82.240 ;
        RECT 104.575 80.840 106.275 82.240 ;
        RECT 106.575 80.840 108.275 82.240 ;
        RECT 108.575 80.840 110.275 82.240 ;
        RECT 110.575 80.840 112.275 82.240 ;
        RECT 112.575 80.840 114.275 82.240 ;
        RECT 114.575 80.840 116.275 82.240 ;
        RECT 116.575 80.840 118.275 82.240 ;
        RECT 118.575 80.840 120.275 82.240 ;
        RECT 120.575 80.840 122.275 82.240 ;
        RECT 122.575 80.840 124.275 82.240 ;
        RECT 124.575 80.840 126.275 82.240 ;
        RECT 126.575 80.840 128.275 82.240 ;
        RECT 128.575 80.840 130.275 82.240 ;
        RECT 130.575 80.840 132.275 82.240 ;
        RECT 132.575 80.840 134.275 82.240 ;
        RECT 134.575 80.840 136.275 82.240 ;
        RECT 136.575 80.840 138.275 82.240 ;
        RECT 138.575 80.840 140.275 82.240 ;
        RECT 140.575 80.840 142.275 82.240 ;
        RECT 142.575 80.840 144.275 82.240 ;
        RECT 144.575 80.840 146.275 82.240 ;
        RECT 146.575 80.840 148.275 82.240 ;
        RECT 148.575 80.840 150.275 82.240 ;
        RECT 150.575 80.840 152.275 82.240 ;
        RECT 152.575 80.840 154.275 82.240 ;
        RECT 6.840 78.990 8.540 80.390 ;
        RECT 8.840 78.990 10.540 80.390 ;
        RECT 10.840 78.990 12.540 80.390 ;
        RECT 12.840 78.990 14.540 80.390 ;
        RECT 14.840 78.990 16.540 80.390 ;
        RECT 16.840 78.990 18.540 80.390 ;
        RECT 18.840 78.990 20.540 80.390 ;
        RECT 20.840 78.990 22.540 80.390 ;
        RECT 22.840 78.990 24.540 80.390 ;
        RECT 24.840 78.990 26.540 80.390 ;
        RECT 26.840 78.990 28.540 80.390 ;
        RECT 28.840 78.990 30.540 80.390 ;
        RECT 30.840 78.990 32.540 80.390 ;
        RECT 32.840 78.990 34.540 80.390 ;
        RECT 34.840 78.990 36.540 80.390 ;
        RECT 36.840 78.990 38.540 80.390 ;
        RECT 38.840 78.990 40.540 80.390 ;
        RECT 40.840 78.990 42.540 80.390 ;
        RECT 42.840 78.990 44.540 80.390 ;
        RECT 44.840 78.990 46.540 80.390 ;
        RECT 46.840 78.990 48.540 80.390 ;
        RECT 48.840 78.990 50.540 80.390 ;
        RECT 50.840 78.990 52.540 80.390 ;
        RECT 52.840 78.990 54.540 80.390 ;
        RECT 54.840 78.990 56.540 80.390 ;
        RECT 56.840 78.990 58.540 80.390 ;
        RECT 58.840 78.990 60.540 80.390 ;
        RECT 60.840 78.990 62.540 80.390 ;
        RECT 62.840 78.990 64.540 80.390 ;
        RECT 64.840 78.990 66.540 80.390 ;
        RECT 66.840 78.990 68.540 80.390 ;
        RECT 68.840 78.990 70.540 80.390 ;
        RECT 70.840 78.990 72.540 80.390 ;
        RECT 72.840 78.990 74.540 80.390 ;
        RECT 86.575 78.990 88.275 80.390 ;
        RECT 88.575 78.990 90.275 80.390 ;
        RECT 90.575 78.990 92.275 80.390 ;
        RECT 92.575 78.990 94.275 80.390 ;
        RECT 94.575 78.990 96.275 80.390 ;
        RECT 96.575 78.990 98.275 80.390 ;
        RECT 98.575 78.990 100.275 80.390 ;
        RECT 100.575 78.990 102.275 80.390 ;
        RECT 102.575 78.990 104.275 80.390 ;
        RECT 104.575 78.990 106.275 80.390 ;
        RECT 106.575 78.990 108.275 80.390 ;
        RECT 108.575 78.990 110.275 80.390 ;
        RECT 110.575 78.990 112.275 80.390 ;
        RECT 112.575 78.990 114.275 80.390 ;
        RECT 114.575 78.990 116.275 80.390 ;
        RECT 116.575 78.990 118.275 80.390 ;
        RECT 118.575 78.990 120.275 80.390 ;
        RECT 120.575 78.990 122.275 80.390 ;
        RECT 122.575 78.990 124.275 80.390 ;
        RECT 124.575 78.990 126.275 80.390 ;
        RECT 126.575 78.990 128.275 80.390 ;
        RECT 128.575 78.990 130.275 80.390 ;
        RECT 130.575 78.990 132.275 80.390 ;
        RECT 132.575 78.990 134.275 80.390 ;
        RECT 134.575 78.990 136.275 80.390 ;
        RECT 136.575 78.990 138.275 80.390 ;
        RECT 138.575 78.990 140.275 80.390 ;
        RECT 140.575 78.990 142.275 80.390 ;
        RECT 142.575 78.990 144.275 80.390 ;
        RECT 144.575 78.990 146.275 80.390 ;
        RECT 146.575 78.990 148.275 80.390 ;
        RECT 148.575 78.990 150.275 80.390 ;
        RECT 150.575 78.990 152.275 80.390 ;
        RECT 152.575 78.990 154.275 80.390 ;
        RECT 6.840 77.140 8.540 78.540 ;
        RECT 8.840 77.140 10.540 78.540 ;
        RECT 10.840 77.140 12.540 78.540 ;
        RECT 12.840 77.140 14.540 78.540 ;
        RECT 14.840 77.140 16.540 78.540 ;
        RECT 16.840 77.140 18.540 78.540 ;
        RECT 18.840 77.140 20.540 78.540 ;
        RECT 20.840 77.140 22.540 78.540 ;
        RECT 22.840 77.140 24.540 78.540 ;
        RECT 24.840 77.140 26.540 78.540 ;
        RECT 26.840 77.140 28.540 78.540 ;
        RECT 28.840 77.140 30.540 78.540 ;
        RECT 30.840 77.140 32.540 78.540 ;
        RECT 32.840 77.140 34.540 78.540 ;
        RECT 34.840 77.140 36.540 78.540 ;
        RECT 36.840 77.140 38.540 78.540 ;
        RECT 38.840 77.140 40.540 78.540 ;
        RECT 40.840 77.140 42.540 78.540 ;
        RECT 42.840 77.140 44.540 78.540 ;
        RECT 44.840 77.140 46.540 78.540 ;
        RECT 46.840 77.140 48.540 78.540 ;
        RECT 48.840 77.140 50.540 78.540 ;
        RECT 50.840 77.140 52.540 78.540 ;
        RECT 52.840 77.140 54.540 78.540 ;
        RECT 54.840 77.140 56.540 78.540 ;
        RECT 56.840 77.140 58.540 78.540 ;
        RECT 58.840 77.140 60.540 78.540 ;
        RECT 60.840 77.140 62.540 78.540 ;
        RECT 62.840 77.140 64.540 78.540 ;
        RECT 64.840 77.140 66.540 78.540 ;
        RECT 66.840 77.140 68.540 78.540 ;
        RECT 68.840 77.140 70.540 78.540 ;
        RECT 70.840 77.140 72.540 78.540 ;
        RECT 72.840 77.140 74.540 78.540 ;
        RECT 86.575 77.140 88.275 78.540 ;
        RECT 88.575 77.140 90.275 78.540 ;
        RECT 90.575 77.140 92.275 78.540 ;
        RECT 92.575 77.140 94.275 78.540 ;
        RECT 94.575 77.140 96.275 78.540 ;
        RECT 96.575 77.140 98.275 78.540 ;
        RECT 98.575 77.140 100.275 78.540 ;
        RECT 100.575 77.140 102.275 78.540 ;
        RECT 102.575 77.140 104.275 78.540 ;
        RECT 104.575 77.140 106.275 78.540 ;
        RECT 106.575 77.140 108.275 78.540 ;
        RECT 108.575 77.140 110.275 78.540 ;
        RECT 110.575 77.140 112.275 78.540 ;
        RECT 112.575 77.140 114.275 78.540 ;
        RECT 114.575 77.140 116.275 78.540 ;
        RECT 116.575 77.140 118.275 78.540 ;
        RECT 118.575 77.140 120.275 78.540 ;
        RECT 120.575 77.140 122.275 78.540 ;
        RECT 122.575 77.140 124.275 78.540 ;
        RECT 124.575 77.140 126.275 78.540 ;
        RECT 126.575 77.140 128.275 78.540 ;
        RECT 128.575 77.140 130.275 78.540 ;
        RECT 130.575 77.140 132.275 78.540 ;
        RECT 132.575 77.140 134.275 78.540 ;
        RECT 134.575 77.140 136.275 78.540 ;
        RECT 136.575 77.140 138.275 78.540 ;
        RECT 138.575 77.140 140.275 78.540 ;
        RECT 140.575 77.140 142.275 78.540 ;
        RECT 142.575 77.140 144.275 78.540 ;
        RECT 144.575 77.140 146.275 78.540 ;
        RECT 146.575 77.140 148.275 78.540 ;
        RECT 148.575 77.140 150.275 78.540 ;
        RECT 150.575 77.140 152.275 78.540 ;
        RECT 152.575 77.140 154.275 78.540 ;
        RECT 6.840 75.290 8.540 76.690 ;
        RECT 8.840 75.290 10.540 76.690 ;
        RECT 10.840 75.290 12.540 76.690 ;
        RECT 12.840 75.290 14.540 76.690 ;
        RECT 14.840 75.290 16.540 76.690 ;
        RECT 16.840 75.290 18.540 76.690 ;
        RECT 18.840 75.290 20.540 76.690 ;
        RECT 20.840 75.290 22.540 76.690 ;
        RECT 22.840 75.290 24.540 76.690 ;
        RECT 24.840 75.290 26.540 76.690 ;
        RECT 26.840 75.290 28.540 76.690 ;
        RECT 28.840 75.290 30.540 76.690 ;
        RECT 30.840 75.290 32.540 76.690 ;
        RECT 32.840 75.290 34.540 76.690 ;
        RECT 34.840 75.290 36.540 76.690 ;
        RECT 36.840 75.290 38.540 76.690 ;
        RECT 38.840 75.290 40.540 76.690 ;
        RECT 40.840 75.290 42.540 76.690 ;
        RECT 42.840 75.290 44.540 76.690 ;
        RECT 44.840 75.290 46.540 76.690 ;
        RECT 46.840 75.290 48.540 76.690 ;
        RECT 48.840 75.290 50.540 76.690 ;
        RECT 50.840 75.290 52.540 76.690 ;
        RECT 52.840 75.290 54.540 76.690 ;
        RECT 54.840 75.290 56.540 76.690 ;
        RECT 56.840 75.290 58.540 76.690 ;
        RECT 58.840 75.290 60.540 76.690 ;
        RECT 60.840 75.290 62.540 76.690 ;
        RECT 62.840 75.290 64.540 76.690 ;
        RECT 64.840 75.290 66.540 76.690 ;
        RECT 66.840 75.290 68.540 76.690 ;
        RECT 68.840 75.290 70.540 76.690 ;
        RECT 70.840 75.290 72.540 76.690 ;
        RECT 72.840 75.290 74.540 76.690 ;
        RECT 86.575 75.290 88.275 76.690 ;
        RECT 88.575 75.290 90.275 76.690 ;
        RECT 90.575 75.290 92.275 76.690 ;
        RECT 92.575 75.290 94.275 76.690 ;
        RECT 94.575 75.290 96.275 76.690 ;
        RECT 96.575 75.290 98.275 76.690 ;
        RECT 98.575 75.290 100.275 76.690 ;
        RECT 100.575 75.290 102.275 76.690 ;
        RECT 102.575 75.290 104.275 76.690 ;
        RECT 104.575 75.290 106.275 76.690 ;
        RECT 106.575 75.290 108.275 76.690 ;
        RECT 108.575 75.290 110.275 76.690 ;
        RECT 110.575 75.290 112.275 76.690 ;
        RECT 112.575 75.290 114.275 76.690 ;
        RECT 114.575 75.290 116.275 76.690 ;
        RECT 116.575 75.290 118.275 76.690 ;
        RECT 118.575 75.290 120.275 76.690 ;
        RECT 120.575 75.290 122.275 76.690 ;
        RECT 122.575 75.290 124.275 76.690 ;
        RECT 124.575 75.290 126.275 76.690 ;
        RECT 126.575 75.290 128.275 76.690 ;
        RECT 128.575 75.290 130.275 76.690 ;
        RECT 130.575 75.290 132.275 76.690 ;
        RECT 132.575 75.290 134.275 76.690 ;
        RECT 134.575 75.290 136.275 76.690 ;
        RECT 136.575 75.290 138.275 76.690 ;
        RECT 138.575 75.290 140.275 76.690 ;
        RECT 140.575 75.290 142.275 76.690 ;
        RECT 142.575 75.290 144.275 76.690 ;
        RECT 144.575 75.290 146.275 76.690 ;
        RECT 146.575 75.290 148.275 76.690 ;
        RECT 148.575 75.290 150.275 76.690 ;
        RECT 150.575 75.290 152.275 76.690 ;
        RECT 152.575 75.290 154.275 76.690 ;
        RECT 6.840 73.440 8.540 74.840 ;
        RECT 8.840 73.440 10.540 74.840 ;
        RECT 10.840 73.440 12.540 74.840 ;
        RECT 12.840 73.440 14.540 74.840 ;
        RECT 14.840 73.440 16.540 74.840 ;
        RECT 16.840 73.440 18.540 74.840 ;
        RECT 18.840 73.440 20.540 74.840 ;
        RECT 20.840 73.440 22.540 74.840 ;
        RECT 22.840 73.440 24.540 74.840 ;
        RECT 24.840 73.440 26.540 74.840 ;
        RECT 26.840 73.440 28.540 74.840 ;
        RECT 28.840 73.440 30.540 74.840 ;
        RECT 30.840 73.440 32.540 74.840 ;
        RECT 32.840 73.440 34.540 74.840 ;
        RECT 34.840 73.440 36.540 74.840 ;
        RECT 36.840 73.440 38.540 74.840 ;
        RECT 38.840 73.440 40.540 74.840 ;
        RECT 40.840 73.440 42.540 74.840 ;
        RECT 42.840 73.440 44.540 74.840 ;
        RECT 44.840 73.440 46.540 74.840 ;
        RECT 46.840 73.440 48.540 74.840 ;
        RECT 48.840 73.440 50.540 74.840 ;
        RECT 50.840 73.440 52.540 74.840 ;
        RECT 52.840 73.440 54.540 74.840 ;
        RECT 54.840 73.440 56.540 74.840 ;
        RECT 56.840 73.440 58.540 74.840 ;
        RECT 58.840 73.440 60.540 74.840 ;
        RECT 60.840 73.440 62.540 74.840 ;
        RECT 62.840 73.440 64.540 74.840 ;
        RECT 64.840 73.440 66.540 74.840 ;
        RECT 66.840 73.440 68.540 74.840 ;
        RECT 68.840 73.440 70.540 74.840 ;
        RECT 70.840 73.440 72.540 74.840 ;
        RECT 72.840 73.440 74.540 74.840 ;
        RECT 86.575 73.440 88.275 74.840 ;
        RECT 88.575 73.440 90.275 74.840 ;
        RECT 90.575 73.440 92.275 74.840 ;
        RECT 92.575 73.440 94.275 74.840 ;
        RECT 94.575 73.440 96.275 74.840 ;
        RECT 96.575 73.440 98.275 74.840 ;
        RECT 98.575 73.440 100.275 74.840 ;
        RECT 100.575 73.440 102.275 74.840 ;
        RECT 102.575 73.440 104.275 74.840 ;
        RECT 104.575 73.440 106.275 74.840 ;
        RECT 106.575 73.440 108.275 74.840 ;
        RECT 108.575 73.440 110.275 74.840 ;
        RECT 110.575 73.440 112.275 74.840 ;
        RECT 112.575 73.440 114.275 74.840 ;
        RECT 114.575 73.440 116.275 74.840 ;
        RECT 116.575 73.440 118.275 74.840 ;
        RECT 118.575 73.440 120.275 74.840 ;
        RECT 120.575 73.440 122.275 74.840 ;
        RECT 122.575 73.440 124.275 74.840 ;
        RECT 124.575 73.440 126.275 74.840 ;
        RECT 126.575 73.440 128.275 74.840 ;
        RECT 128.575 73.440 130.275 74.840 ;
        RECT 130.575 73.440 132.275 74.840 ;
        RECT 132.575 73.440 134.275 74.840 ;
        RECT 134.575 73.440 136.275 74.840 ;
        RECT 136.575 73.440 138.275 74.840 ;
        RECT 138.575 73.440 140.275 74.840 ;
        RECT 140.575 73.440 142.275 74.840 ;
        RECT 142.575 73.440 144.275 74.840 ;
        RECT 144.575 73.440 146.275 74.840 ;
        RECT 146.575 73.440 148.275 74.840 ;
        RECT 148.575 73.440 150.275 74.840 ;
        RECT 150.575 73.440 152.275 74.840 ;
        RECT 152.575 73.440 154.275 74.840 ;
        RECT 6.840 71.590 8.540 72.990 ;
        RECT 8.840 71.590 10.540 72.990 ;
        RECT 10.840 71.590 12.540 72.990 ;
        RECT 12.840 71.590 14.540 72.990 ;
        RECT 14.840 71.590 16.540 72.990 ;
        RECT 16.840 71.590 18.540 72.990 ;
        RECT 18.840 71.590 20.540 72.990 ;
        RECT 20.840 71.590 22.540 72.990 ;
        RECT 22.840 71.590 24.540 72.990 ;
        RECT 24.840 71.590 26.540 72.990 ;
        RECT 26.840 71.590 28.540 72.990 ;
        RECT 28.840 71.590 30.540 72.990 ;
        RECT 30.840 71.590 32.540 72.990 ;
        RECT 32.840 71.590 34.540 72.990 ;
        RECT 34.840 71.590 36.540 72.990 ;
        RECT 36.840 71.590 38.540 72.990 ;
        RECT 38.840 71.590 40.540 72.990 ;
        RECT 40.840 71.590 42.540 72.990 ;
        RECT 42.840 71.590 44.540 72.990 ;
        RECT 44.840 71.590 46.540 72.990 ;
        RECT 46.840 71.590 48.540 72.990 ;
        RECT 48.840 71.590 50.540 72.990 ;
        RECT 50.840 71.590 52.540 72.990 ;
        RECT 52.840 71.590 54.540 72.990 ;
        RECT 54.840 71.590 56.540 72.990 ;
        RECT 56.840 71.590 58.540 72.990 ;
        RECT 58.840 71.590 60.540 72.990 ;
        RECT 60.840 71.590 62.540 72.990 ;
        RECT 62.840 71.590 64.540 72.990 ;
        RECT 64.840 71.590 66.540 72.990 ;
        RECT 66.840 71.590 68.540 72.990 ;
        RECT 68.840 71.590 70.540 72.990 ;
        RECT 70.840 71.590 72.540 72.990 ;
        RECT 72.840 71.590 74.540 72.990 ;
        RECT 86.575 71.590 88.275 72.990 ;
        RECT 88.575 71.590 90.275 72.990 ;
        RECT 90.575 71.590 92.275 72.990 ;
        RECT 92.575 71.590 94.275 72.990 ;
        RECT 94.575 71.590 96.275 72.990 ;
        RECT 96.575 71.590 98.275 72.990 ;
        RECT 98.575 71.590 100.275 72.990 ;
        RECT 100.575 71.590 102.275 72.990 ;
        RECT 102.575 71.590 104.275 72.990 ;
        RECT 104.575 71.590 106.275 72.990 ;
        RECT 106.575 71.590 108.275 72.990 ;
        RECT 108.575 71.590 110.275 72.990 ;
        RECT 110.575 71.590 112.275 72.990 ;
        RECT 112.575 71.590 114.275 72.990 ;
        RECT 114.575 71.590 116.275 72.990 ;
        RECT 116.575 71.590 118.275 72.990 ;
        RECT 118.575 71.590 120.275 72.990 ;
        RECT 120.575 71.590 122.275 72.990 ;
        RECT 122.575 71.590 124.275 72.990 ;
        RECT 124.575 71.590 126.275 72.990 ;
        RECT 126.575 71.590 128.275 72.990 ;
        RECT 128.575 71.590 130.275 72.990 ;
        RECT 130.575 71.590 132.275 72.990 ;
        RECT 132.575 71.590 134.275 72.990 ;
        RECT 134.575 71.590 136.275 72.990 ;
        RECT 136.575 71.590 138.275 72.990 ;
        RECT 138.575 71.590 140.275 72.990 ;
        RECT 140.575 71.590 142.275 72.990 ;
        RECT 142.575 71.590 144.275 72.990 ;
        RECT 144.575 71.590 146.275 72.990 ;
        RECT 146.575 71.590 148.275 72.990 ;
        RECT 148.575 71.590 150.275 72.990 ;
        RECT 150.575 71.590 152.275 72.990 ;
        RECT 152.575 71.590 154.275 72.990 ;
        RECT 6.840 69.740 8.540 71.140 ;
        RECT 8.840 69.740 10.540 71.140 ;
        RECT 10.840 69.740 12.540 71.140 ;
        RECT 12.840 69.740 14.540 71.140 ;
        RECT 14.840 69.740 16.540 71.140 ;
        RECT 16.840 69.740 18.540 71.140 ;
        RECT 18.840 69.740 20.540 71.140 ;
        RECT 20.840 69.740 22.540 71.140 ;
        RECT 22.840 69.740 24.540 71.140 ;
        RECT 24.840 69.740 26.540 71.140 ;
        RECT 26.840 69.740 28.540 71.140 ;
        RECT 28.840 69.740 30.540 71.140 ;
        RECT 30.840 69.740 32.540 71.140 ;
        RECT 32.840 69.740 34.540 71.140 ;
        RECT 34.840 69.740 36.540 71.140 ;
        RECT 36.840 69.740 38.540 71.140 ;
        RECT 38.840 69.740 40.540 71.140 ;
        RECT 40.840 69.740 42.540 71.140 ;
        RECT 42.840 69.740 44.540 71.140 ;
        RECT 44.840 69.740 46.540 71.140 ;
        RECT 46.840 69.740 48.540 71.140 ;
        RECT 48.840 69.740 50.540 71.140 ;
        RECT 50.840 69.740 52.540 71.140 ;
        RECT 52.840 69.740 54.540 71.140 ;
        RECT 54.840 69.740 56.540 71.140 ;
        RECT 56.840 69.740 58.540 71.140 ;
        RECT 58.840 69.740 60.540 71.140 ;
        RECT 60.840 69.740 62.540 71.140 ;
        RECT 62.840 69.740 64.540 71.140 ;
        RECT 64.840 69.740 66.540 71.140 ;
        RECT 66.840 69.740 68.540 71.140 ;
        RECT 68.840 69.740 70.540 71.140 ;
        RECT 70.840 69.740 72.540 71.140 ;
        RECT 72.840 69.740 74.540 71.140 ;
        RECT 86.575 69.740 88.275 71.140 ;
        RECT 88.575 69.740 90.275 71.140 ;
        RECT 90.575 69.740 92.275 71.140 ;
        RECT 92.575 69.740 94.275 71.140 ;
        RECT 94.575 69.740 96.275 71.140 ;
        RECT 96.575 69.740 98.275 71.140 ;
        RECT 98.575 69.740 100.275 71.140 ;
        RECT 100.575 69.740 102.275 71.140 ;
        RECT 102.575 69.740 104.275 71.140 ;
        RECT 104.575 69.740 106.275 71.140 ;
        RECT 106.575 69.740 108.275 71.140 ;
        RECT 108.575 69.740 110.275 71.140 ;
        RECT 110.575 69.740 112.275 71.140 ;
        RECT 112.575 69.740 114.275 71.140 ;
        RECT 114.575 69.740 116.275 71.140 ;
        RECT 116.575 69.740 118.275 71.140 ;
        RECT 118.575 69.740 120.275 71.140 ;
        RECT 120.575 69.740 122.275 71.140 ;
        RECT 122.575 69.740 124.275 71.140 ;
        RECT 124.575 69.740 126.275 71.140 ;
        RECT 126.575 69.740 128.275 71.140 ;
        RECT 128.575 69.740 130.275 71.140 ;
        RECT 130.575 69.740 132.275 71.140 ;
        RECT 132.575 69.740 134.275 71.140 ;
        RECT 134.575 69.740 136.275 71.140 ;
        RECT 136.575 69.740 138.275 71.140 ;
        RECT 138.575 69.740 140.275 71.140 ;
        RECT 140.575 69.740 142.275 71.140 ;
        RECT 142.575 69.740 144.275 71.140 ;
        RECT 144.575 69.740 146.275 71.140 ;
        RECT 146.575 69.740 148.275 71.140 ;
        RECT 148.575 69.740 150.275 71.140 ;
        RECT 150.575 69.740 152.275 71.140 ;
        RECT 152.575 69.740 154.275 71.140 ;
        RECT 6.840 67.890 8.540 69.290 ;
        RECT 8.840 67.890 10.540 69.290 ;
        RECT 10.840 67.890 12.540 69.290 ;
        RECT 12.840 67.890 14.540 69.290 ;
        RECT 14.840 67.890 16.540 69.290 ;
        RECT 16.840 67.890 18.540 69.290 ;
        RECT 18.840 67.890 20.540 69.290 ;
        RECT 20.840 67.890 22.540 69.290 ;
        RECT 22.840 67.890 24.540 69.290 ;
        RECT 24.840 67.890 26.540 69.290 ;
        RECT 26.840 67.890 28.540 69.290 ;
        RECT 28.840 67.890 30.540 69.290 ;
        RECT 30.840 67.890 32.540 69.290 ;
        RECT 32.840 67.890 34.540 69.290 ;
        RECT 34.840 67.890 36.540 69.290 ;
        RECT 36.840 67.890 38.540 69.290 ;
        RECT 38.840 67.890 40.540 69.290 ;
        RECT 40.840 67.890 42.540 69.290 ;
        RECT 42.840 67.890 44.540 69.290 ;
        RECT 44.840 67.890 46.540 69.290 ;
        RECT 46.840 67.890 48.540 69.290 ;
        RECT 48.840 67.890 50.540 69.290 ;
        RECT 50.840 67.890 52.540 69.290 ;
        RECT 52.840 67.890 54.540 69.290 ;
        RECT 54.840 67.890 56.540 69.290 ;
        RECT 56.840 67.890 58.540 69.290 ;
        RECT 58.840 67.890 60.540 69.290 ;
        RECT 60.840 67.890 62.540 69.290 ;
        RECT 62.840 67.890 64.540 69.290 ;
        RECT 64.840 67.890 66.540 69.290 ;
        RECT 66.840 67.890 68.540 69.290 ;
        RECT 68.840 67.890 70.540 69.290 ;
        RECT 70.840 67.890 72.540 69.290 ;
        RECT 72.840 67.890 74.540 69.290 ;
        RECT 86.575 67.890 88.275 69.290 ;
        RECT 88.575 67.890 90.275 69.290 ;
        RECT 90.575 67.890 92.275 69.290 ;
        RECT 92.575 67.890 94.275 69.290 ;
        RECT 94.575 67.890 96.275 69.290 ;
        RECT 96.575 67.890 98.275 69.290 ;
        RECT 98.575 67.890 100.275 69.290 ;
        RECT 100.575 67.890 102.275 69.290 ;
        RECT 102.575 67.890 104.275 69.290 ;
        RECT 104.575 67.890 106.275 69.290 ;
        RECT 106.575 67.890 108.275 69.290 ;
        RECT 108.575 67.890 110.275 69.290 ;
        RECT 110.575 67.890 112.275 69.290 ;
        RECT 112.575 67.890 114.275 69.290 ;
        RECT 114.575 67.890 116.275 69.290 ;
        RECT 116.575 67.890 118.275 69.290 ;
        RECT 118.575 67.890 120.275 69.290 ;
        RECT 120.575 67.890 122.275 69.290 ;
        RECT 122.575 67.890 124.275 69.290 ;
        RECT 124.575 67.890 126.275 69.290 ;
        RECT 126.575 67.890 128.275 69.290 ;
        RECT 128.575 67.890 130.275 69.290 ;
        RECT 130.575 67.890 132.275 69.290 ;
        RECT 132.575 67.890 134.275 69.290 ;
        RECT 134.575 67.890 136.275 69.290 ;
        RECT 136.575 67.890 138.275 69.290 ;
        RECT 138.575 67.890 140.275 69.290 ;
        RECT 140.575 67.890 142.275 69.290 ;
        RECT 142.575 67.890 144.275 69.290 ;
        RECT 144.575 67.890 146.275 69.290 ;
        RECT 146.575 67.890 148.275 69.290 ;
        RECT 148.575 67.890 150.275 69.290 ;
        RECT 150.575 67.890 152.275 69.290 ;
        RECT 152.575 67.890 154.275 69.290 ;
        RECT 6.840 66.040 8.540 67.440 ;
        RECT 8.840 66.040 10.540 67.440 ;
        RECT 10.840 66.040 12.540 67.440 ;
        RECT 12.840 66.040 14.540 67.440 ;
        RECT 14.840 66.040 16.540 67.440 ;
        RECT 16.840 66.040 18.540 67.440 ;
        RECT 18.840 66.040 20.540 67.440 ;
        RECT 20.840 66.040 22.540 67.440 ;
        RECT 22.840 66.040 24.540 67.440 ;
        RECT 24.840 66.040 26.540 67.440 ;
        RECT 26.840 66.040 28.540 67.440 ;
        RECT 28.840 66.040 30.540 67.440 ;
        RECT 30.840 66.040 32.540 67.440 ;
        RECT 32.840 66.040 34.540 67.440 ;
        RECT 34.840 66.040 36.540 67.440 ;
        RECT 36.840 66.040 38.540 67.440 ;
        RECT 38.840 66.040 40.540 67.440 ;
        RECT 40.840 66.040 42.540 67.440 ;
        RECT 42.840 66.040 44.540 67.440 ;
        RECT 44.840 66.040 46.540 67.440 ;
        RECT 46.840 66.040 48.540 67.440 ;
        RECT 48.840 66.040 50.540 67.440 ;
        RECT 50.840 66.040 52.540 67.440 ;
        RECT 52.840 66.040 54.540 67.440 ;
        RECT 54.840 66.040 56.540 67.440 ;
        RECT 56.840 66.040 58.540 67.440 ;
        RECT 58.840 66.040 60.540 67.440 ;
        RECT 60.840 66.040 62.540 67.440 ;
        RECT 62.840 66.040 64.540 67.440 ;
        RECT 64.840 66.040 66.540 67.440 ;
        RECT 66.840 66.040 68.540 67.440 ;
        RECT 68.840 66.040 70.540 67.440 ;
        RECT 70.840 66.040 72.540 67.440 ;
        RECT 72.840 66.040 74.540 67.440 ;
        RECT 86.575 66.040 88.275 67.440 ;
        RECT 88.575 66.040 90.275 67.440 ;
        RECT 90.575 66.040 92.275 67.440 ;
        RECT 92.575 66.040 94.275 67.440 ;
        RECT 94.575 66.040 96.275 67.440 ;
        RECT 96.575 66.040 98.275 67.440 ;
        RECT 98.575 66.040 100.275 67.440 ;
        RECT 100.575 66.040 102.275 67.440 ;
        RECT 102.575 66.040 104.275 67.440 ;
        RECT 104.575 66.040 106.275 67.440 ;
        RECT 106.575 66.040 108.275 67.440 ;
        RECT 108.575 66.040 110.275 67.440 ;
        RECT 110.575 66.040 112.275 67.440 ;
        RECT 112.575 66.040 114.275 67.440 ;
        RECT 114.575 66.040 116.275 67.440 ;
        RECT 116.575 66.040 118.275 67.440 ;
        RECT 118.575 66.040 120.275 67.440 ;
        RECT 120.575 66.040 122.275 67.440 ;
        RECT 122.575 66.040 124.275 67.440 ;
        RECT 124.575 66.040 126.275 67.440 ;
        RECT 126.575 66.040 128.275 67.440 ;
        RECT 128.575 66.040 130.275 67.440 ;
        RECT 130.575 66.040 132.275 67.440 ;
        RECT 132.575 66.040 134.275 67.440 ;
        RECT 134.575 66.040 136.275 67.440 ;
        RECT 136.575 66.040 138.275 67.440 ;
        RECT 138.575 66.040 140.275 67.440 ;
        RECT 140.575 66.040 142.275 67.440 ;
        RECT 142.575 66.040 144.275 67.440 ;
        RECT 144.575 66.040 146.275 67.440 ;
        RECT 146.575 66.040 148.275 67.440 ;
        RECT 148.575 66.040 150.275 67.440 ;
        RECT 150.575 66.040 152.275 67.440 ;
        RECT 152.575 66.040 154.275 67.440 ;
        RECT 6.840 64.190 8.540 65.590 ;
        RECT 8.840 64.190 10.540 65.590 ;
        RECT 10.840 64.190 12.540 65.590 ;
        RECT 12.840 64.190 14.540 65.590 ;
        RECT 14.840 64.190 16.540 65.590 ;
        RECT 16.840 64.190 18.540 65.590 ;
        RECT 18.840 64.190 20.540 65.590 ;
        RECT 20.840 64.190 22.540 65.590 ;
        RECT 22.840 64.190 24.540 65.590 ;
        RECT 24.840 64.190 26.540 65.590 ;
        RECT 26.840 64.190 28.540 65.590 ;
        RECT 28.840 64.190 30.540 65.590 ;
        RECT 30.840 64.190 32.540 65.590 ;
        RECT 32.840 64.190 34.540 65.590 ;
        RECT 34.840 64.190 36.540 65.590 ;
        RECT 36.840 64.190 38.540 65.590 ;
        RECT 38.840 64.190 40.540 65.590 ;
        RECT 40.840 64.190 42.540 65.590 ;
        RECT 42.840 64.190 44.540 65.590 ;
        RECT 44.840 64.190 46.540 65.590 ;
        RECT 46.840 64.190 48.540 65.590 ;
        RECT 48.840 64.190 50.540 65.590 ;
        RECT 50.840 64.190 52.540 65.590 ;
        RECT 52.840 64.190 54.540 65.590 ;
        RECT 54.840 64.190 56.540 65.590 ;
        RECT 56.840 64.190 58.540 65.590 ;
        RECT 58.840 64.190 60.540 65.590 ;
        RECT 60.840 64.190 62.540 65.590 ;
        RECT 62.840 64.190 64.540 65.590 ;
        RECT 64.840 64.190 66.540 65.590 ;
        RECT 66.840 64.190 68.540 65.590 ;
        RECT 68.840 64.190 70.540 65.590 ;
        RECT 70.840 64.190 72.540 65.590 ;
        RECT 72.840 64.190 74.540 65.590 ;
        RECT 86.575 64.190 88.275 65.590 ;
        RECT 88.575 64.190 90.275 65.590 ;
        RECT 90.575 64.190 92.275 65.590 ;
        RECT 92.575 64.190 94.275 65.590 ;
        RECT 94.575 64.190 96.275 65.590 ;
        RECT 96.575 64.190 98.275 65.590 ;
        RECT 98.575 64.190 100.275 65.590 ;
        RECT 100.575 64.190 102.275 65.590 ;
        RECT 102.575 64.190 104.275 65.590 ;
        RECT 104.575 64.190 106.275 65.590 ;
        RECT 106.575 64.190 108.275 65.590 ;
        RECT 108.575 64.190 110.275 65.590 ;
        RECT 110.575 64.190 112.275 65.590 ;
        RECT 112.575 64.190 114.275 65.590 ;
        RECT 114.575 64.190 116.275 65.590 ;
        RECT 116.575 64.190 118.275 65.590 ;
        RECT 118.575 64.190 120.275 65.590 ;
        RECT 120.575 64.190 122.275 65.590 ;
        RECT 122.575 64.190 124.275 65.590 ;
        RECT 124.575 64.190 126.275 65.590 ;
        RECT 126.575 64.190 128.275 65.590 ;
        RECT 128.575 64.190 130.275 65.590 ;
        RECT 130.575 64.190 132.275 65.590 ;
        RECT 132.575 64.190 134.275 65.590 ;
        RECT 134.575 64.190 136.275 65.590 ;
        RECT 136.575 64.190 138.275 65.590 ;
        RECT 138.575 64.190 140.275 65.590 ;
        RECT 140.575 64.190 142.275 65.590 ;
        RECT 142.575 64.190 144.275 65.590 ;
        RECT 144.575 64.190 146.275 65.590 ;
        RECT 146.575 64.190 148.275 65.590 ;
        RECT 148.575 64.190 150.275 65.590 ;
        RECT 150.575 64.190 152.275 65.590 ;
        RECT 152.575 64.190 154.275 65.590 ;
        RECT 6.840 62.340 8.540 63.740 ;
        RECT 8.840 62.340 10.540 63.740 ;
        RECT 10.840 62.340 12.540 63.740 ;
        RECT 12.840 62.340 14.540 63.740 ;
        RECT 14.840 62.340 16.540 63.740 ;
        RECT 16.840 62.340 18.540 63.740 ;
        RECT 18.840 62.340 20.540 63.740 ;
        RECT 20.840 62.340 22.540 63.740 ;
        RECT 22.840 62.340 24.540 63.740 ;
        RECT 24.840 62.340 26.540 63.740 ;
        RECT 26.840 62.340 28.540 63.740 ;
        RECT 28.840 62.340 30.540 63.740 ;
        RECT 30.840 62.340 32.540 63.740 ;
        RECT 32.840 62.340 34.540 63.740 ;
        RECT 34.840 62.340 36.540 63.740 ;
        RECT 36.840 62.340 38.540 63.740 ;
        RECT 38.840 62.340 40.540 63.740 ;
        RECT 40.840 62.340 42.540 63.740 ;
        RECT 42.840 62.340 44.540 63.740 ;
        RECT 44.840 62.340 46.540 63.740 ;
        RECT 46.840 62.340 48.540 63.740 ;
        RECT 48.840 62.340 50.540 63.740 ;
        RECT 50.840 62.340 52.540 63.740 ;
        RECT 52.840 62.340 54.540 63.740 ;
        RECT 54.840 62.340 56.540 63.740 ;
        RECT 56.840 62.340 58.540 63.740 ;
        RECT 58.840 62.340 60.540 63.740 ;
        RECT 60.840 62.340 62.540 63.740 ;
        RECT 62.840 62.340 64.540 63.740 ;
        RECT 64.840 62.340 66.540 63.740 ;
        RECT 66.840 62.340 68.540 63.740 ;
        RECT 68.840 62.340 70.540 63.740 ;
        RECT 70.840 62.340 72.540 63.740 ;
        RECT 72.840 62.340 74.540 63.740 ;
        RECT 86.575 62.340 88.275 63.740 ;
        RECT 88.575 62.340 90.275 63.740 ;
        RECT 90.575 62.340 92.275 63.740 ;
        RECT 92.575 62.340 94.275 63.740 ;
        RECT 94.575 62.340 96.275 63.740 ;
        RECT 96.575 62.340 98.275 63.740 ;
        RECT 98.575 62.340 100.275 63.740 ;
        RECT 100.575 62.340 102.275 63.740 ;
        RECT 102.575 62.340 104.275 63.740 ;
        RECT 104.575 62.340 106.275 63.740 ;
        RECT 106.575 62.340 108.275 63.740 ;
        RECT 108.575 62.340 110.275 63.740 ;
        RECT 110.575 62.340 112.275 63.740 ;
        RECT 112.575 62.340 114.275 63.740 ;
        RECT 114.575 62.340 116.275 63.740 ;
        RECT 116.575 62.340 118.275 63.740 ;
        RECT 118.575 62.340 120.275 63.740 ;
        RECT 120.575 62.340 122.275 63.740 ;
        RECT 122.575 62.340 124.275 63.740 ;
        RECT 124.575 62.340 126.275 63.740 ;
        RECT 126.575 62.340 128.275 63.740 ;
        RECT 128.575 62.340 130.275 63.740 ;
        RECT 130.575 62.340 132.275 63.740 ;
        RECT 132.575 62.340 134.275 63.740 ;
        RECT 134.575 62.340 136.275 63.740 ;
        RECT 136.575 62.340 138.275 63.740 ;
        RECT 138.575 62.340 140.275 63.740 ;
        RECT 140.575 62.340 142.275 63.740 ;
        RECT 142.575 62.340 144.275 63.740 ;
        RECT 144.575 62.340 146.275 63.740 ;
        RECT 146.575 62.340 148.275 63.740 ;
        RECT 148.575 62.340 150.275 63.740 ;
        RECT 150.575 62.340 152.275 63.740 ;
        RECT 152.575 62.340 154.275 63.740 ;
        RECT 6.840 60.490 8.540 61.890 ;
        RECT 8.840 60.490 10.540 61.890 ;
        RECT 10.840 60.490 12.540 61.890 ;
        RECT 12.840 60.490 14.540 61.890 ;
        RECT 14.840 60.490 16.540 61.890 ;
        RECT 16.840 60.490 18.540 61.890 ;
        RECT 18.840 60.490 20.540 61.890 ;
        RECT 20.840 60.490 22.540 61.890 ;
        RECT 22.840 60.490 24.540 61.890 ;
        RECT 24.840 60.490 26.540 61.890 ;
        RECT 26.840 60.490 28.540 61.890 ;
        RECT 28.840 60.490 30.540 61.890 ;
        RECT 30.840 60.490 32.540 61.890 ;
        RECT 32.840 60.490 34.540 61.890 ;
        RECT 34.840 60.490 36.540 61.890 ;
        RECT 36.840 60.490 38.540 61.890 ;
        RECT 38.840 60.490 40.540 61.890 ;
        RECT 40.840 60.490 42.540 61.890 ;
        RECT 42.840 60.490 44.540 61.890 ;
        RECT 44.840 60.490 46.540 61.890 ;
        RECT 46.840 60.490 48.540 61.890 ;
        RECT 48.840 60.490 50.540 61.890 ;
        RECT 50.840 60.490 52.540 61.890 ;
        RECT 52.840 60.490 54.540 61.890 ;
        RECT 54.840 60.490 56.540 61.890 ;
        RECT 56.840 60.490 58.540 61.890 ;
        RECT 58.840 60.490 60.540 61.890 ;
        RECT 60.840 60.490 62.540 61.890 ;
        RECT 62.840 60.490 64.540 61.890 ;
        RECT 64.840 60.490 66.540 61.890 ;
        RECT 66.840 60.490 68.540 61.890 ;
        RECT 68.840 60.490 70.540 61.890 ;
        RECT 70.840 60.490 72.540 61.890 ;
        RECT 72.840 60.490 74.540 61.890 ;
        RECT 86.575 60.490 88.275 61.890 ;
        RECT 88.575 60.490 90.275 61.890 ;
        RECT 90.575 60.490 92.275 61.890 ;
        RECT 92.575 60.490 94.275 61.890 ;
        RECT 94.575 60.490 96.275 61.890 ;
        RECT 96.575 60.490 98.275 61.890 ;
        RECT 98.575 60.490 100.275 61.890 ;
        RECT 100.575 60.490 102.275 61.890 ;
        RECT 102.575 60.490 104.275 61.890 ;
        RECT 104.575 60.490 106.275 61.890 ;
        RECT 106.575 60.490 108.275 61.890 ;
        RECT 108.575 60.490 110.275 61.890 ;
        RECT 110.575 60.490 112.275 61.890 ;
        RECT 112.575 60.490 114.275 61.890 ;
        RECT 114.575 60.490 116.275 61.890 ;
        RECT 116.575 60.490 118.275 61.890 ;
        RECT 118.575 60.490 120.275 61.890 ;
        RECT 120.575 60.490 122.275 61.890 ;
        RECT 122.575 60.490 124.275 61.890 ;
        RECT 124.575 60.490 126.275 61.890 ;
        RECT 126.575 60.490 128.275 61.890 ;
        RECT 128.575 60.490 130.275 61.890 ;
        RECT 130.575 60.490 132.275 61.890 ;
        RECT 132.575 60.490 134.275 61.890 ;
        RECT 134.575 60.490 136.275 61.890 ;
        RECT 136.575 60.490 138.275 61.890 ;
        RECT 138.575 60.490 140.275 61.890 ;
        RECT 140.575 60.490 142.275 61.890 ;
        RECT 142.575 60.490 144.275 61.890 ;
        RECT 144.575 60.490 146.275 61.890 ;
        RECT 146.575 60.490 148.275 61.890 ;
        RECT 148.575 60.490 150.275 61.890 ;
        RECT 150.575 60.490 152.275 61.890 ;
        RECT 152.575 60.490 154.275 61.890 ;
        RECT 6.840 58.640 8.540 60.040 ;
        RECT 8.840 58.640 10.540 60.040 ;
        RECT 10.840 58.640 12.540 60.040 ;
        RECT 12.840 58.640 14.540 60.040 ;
        RECT 14.840 58.640 16.540 60.040 ;
        RECT 16.840 58.640 18.540 60.040 ;
        RECT 18.840 58.640 20.540 60.040 ;
        RECT 20.840 58.640 22.540 60.040 ;
        RECT 22.840 58.640 24.540 60.040 ;
        RECT 24.840 58.640 26.540 60.040 ;
        RECT 26.840 58.640 28.540 60.040 ;
        RECT 28.840 58.640 30.540 60.040 ;
        RECT 30.840 58.640 32.540 60.040 ;
        RECT 32.840 58.640 34.540 60.040 ;
        RECT 34.840 58.640 36.540 60.040 ;
        RECT 36.840 58.640 38.540 60.040 ;
        RECT 38.840 58.640 40.540 60.040 ;
        RECT 40.840 58.640 42.540 60.040 ;
        RECT 42.840 58.640 44.540 60.040 ;
        RECT 44.840 58.640 46.540 60.040 ;
        RECT 46.840 58.640 48.540 60.040 ;
        RECT 48.840 58.640 50.540 60.040 ;
        RECT 50.840 58.640 52.540 60.040 ;
        RECT 52.840 58.640 54.540 60.040 ;
        RECT 54.840 58.640 56.540 60.040 ;
        RECT 56.840 58.640 58.540 60.040 ;
        RECT 58.840 58.640 60.540 60.040 ;
        RECT 60.840 58.640 62.540 60.040 ;
        RECT 62.840 58.640 64.540 60.040 ;
        RECT 64.840 58.640 66.540 60.040 ;
        RECT 66.840 58.640 68.540 60.040 ;
        RECT 68.840 58.640 70.540 60.040 ;
        RECT 70.840 58.640 72.540 60.040 ;
        RECT 72.840 58.640 74.540 60.040 ;
        RECT 86.575 58.640 88.275 60.040 ;
        RECT 88.575 58.640 90.275 60.040 ;
        RECT 90.575 58.640 92.275 60.040 ;
        RECT 92.575 58.640 94.275 60.040 ;
        RECT 94.575 58.640 96.275 60.040 ;
        RECT 96.575 58.640 98.275 60.040 ;
        RECT 98.575 58.640 100.275 60.040 ;
        RECT 100.575 58.640 102.275 60.040 ;
        RECT 102.575 58.640 104.275 60.040 ;
        RECT 104.575 58.640 106.275 60.040 ;
        RECT 106.575 58.640 108.275 60.040 ;
        RECT 108.575 58.640 110.275 60.040 ;
        RECT 110.575 58.640 112.275 60.040 ;
        RECT 112.575 58.640 114.275 60.040 ;
        RECT 114.575 58.640 116.275 60.040 ;
        RECT 116.575 58.640 118.275 60.040 ;
        RECT 118.575 58.640 120.275 60.040 ;
        RECT 120.575 58.640 122.275 60.040 ;
        RECT 122.575 58.640 124.275 60.040 ;
        RECT 124.575 58.640 126.275 60.040 ;
        RECT 126.575 58.640 128.275 60.040 ;
        RECT 128.575 58.640 130.275 60.040 ;
        RECT 130.575 58.640 132.275 60.040 ;
        RECT 132.575 58.640 134.275 60.040 ;
        RECT 134.575 58.640 136.275 60.040 ;
        RECT 136.575 58.640 138.275 60.040 ;
        RECT 138.575 58.640 140.275 60.040 ;
        RECT 140.575 58.640 142.275 60.040 ;
        RECT 142.575 58.640 144.275 60.040 ;
        RECT 144.575 58.640 146.275 60.040 ;
        RECT 146.575 58.640 148.275 60.040 ;
        RECT 148.575 58.640 150.275 60.040 ;
        RECT 150.575 58.640 152.275 60.040 ;
        RECT 152.575 58.640 154.275 60.040 ;
        RECT 6.840 56.790 8.540 58.190 ;
        RECT 8.840 56.790 10.540 58.190 ;
        RECT 10.840 56.790 12.540 58.190 ;
        RECT 12.840 56.790 14.540 58.190 ;
        RECT 14.840 56.790 16.540 58.190 ;
        RECT 16.840 56.790 18.540 58.190 ;
        RECT 18.840 56.790 20.540 58.190 ;
        RECT 20.840 56.790 22.540 58.190 ;
        RECT 22.840 56.790 24.540 58.190 ;
        RECT 24.840 56.790 26.540 58.190 ;
        RECT 26.840 56.790 28.540 58.190 ;
        RECT 28.840 56.790 30.540 58.190 ;
        RECT 30.840 56.790 32.540 58.190 ;
        RECT 32.840 56.790 34.540 58.190 ;
        RECT 34.840 56.790 36.540 58.190 ;
        RECT 36.840 56.790 38.540 58.190 ;
        RECT 38.840 56.790 40.540 58.190 ;
        RECT 40.840 56.790 42.540 58.190 ;
        RECT 42.840 56.790 44.540 58.190 ;
        RECT 44.840 56.790 46.540 58.190 ;
        RECT 46.840 56.790 48.540 58.190 ;
        RECT 48.840 56.790 50.540 58.190 ;
        RECT 50.840 56.790 52.540 58.190 ;
        RECT 52.840 56.790 54.540 58.190 ;
        RECT 54.840 56.790 56.540 58.190 ;
        RECT 56.840 56.790 58.540 58.190 ;
        RECT 58.840 56.790 60.540 58.190 ;
        RECT 60.840 56.790 62.540 58.190 ;
        RECT 62.840 56.790 64.540 58.190 ;
        RECT 64.840 56.790 66.540 58.190 ;
        RECT 66.840 56.790 68.540 58.190 ;
        RECT 68.840 56.790 70.540 58.190 ;
        RECT 70.840 56.790 72.540 58.190 ;
        RECT 72.840 56.790 74.540 58.190 ;
        RECT 86.575 56.790 88.275 58.190 ;
        RECT 88.575 56.790 90.275 58.190 ;
        RECT 90.575 56.790 92.275 58.190 ;
        RECT 92.575 56.790 94.275 58.190 ;
        RECT 94.575 56.790 96.275 58.190 ;
        RECT 96.575 56.790 98.275 58.190 ;
        RECT 98.575 56.790 100.275 58.190 ;
        RECT 100.575 56.790 102.275 58.190 ;
        RECT 102.575 56.790 104.275 58.190 ;
        RECT 104.575 56.790 106.275 58.190 ;
        RECT 106.575 56.790 108.275 58.190 ;
        RECT 108.575 56.790 110.275 58.190 ;
        RECT 110.575 56.790 112.275 58.190 ;
        RECT 112.575 56.790 114.275 58.190 ;
        RECT 114.575 56.790 116.275 58.190 ;
        RECT 116.575 56.790 118.275 58.190 ;
        RECT 118.575 56.790 120.275 58.190 ;
        RECT 120.575 56.790 122.275 58.190 ;
        RECT 122.575 56.790 124.275 58.190 ;
        RECT 124.575 56.790 126.275 58.190 ;
        RECT 126.575 56.790 128.275 58.190 ;
        RECT 128.575 56.790 130.275 58.190 ;
        RECT 130.575 56.790 132.275 58.190 ;
        RECT 132.575 56.790 134.275 58.190 ;
        RECT 134.575 56.790 136.275 58.190 ;
        RECT 136.575 56.790 138.275 58.190 ;
        RECT 138.575 56.790 140.275 58.190 ;
        RECT 140.575 56.790 142.275 58.190 ;
        RECT 142.575 56.790 144.275 58.190 ;
        RECT 144.575 56.790 146.275 58.190 ;
        RECT 146.575 56.790 148.275 58.190 ;
        RECT 148.575 56.790 150.275 58.190 ;
        RECT 150.575 56.790 152.275 58.190 ;
        RECT 152.575 56.790 154.275 58.190 ;
        RECT 6.840 54.940 8.540 56.340 ;
        RECT 8.840 54.940 10.540 56.340 ;
        RECT 10.840 54.940 12.540 56.340 ;
        RECT 12.840 54.940 14.540 56.340 ;
        RECT 14.840 54.940 16.540 56.340 ;
        RECT 16.840 54.940 18.540 56.340 ;
        RECT 18.840 54.940 20.540 56.340 ;
        RECT 20.840 54.940 22.540 56.340 ;
        RECT 22.840 54.940 24.540 56.340 ;
        RECT 24.840 54.940 26.540 56.340 ;
        RECT 26.840 54.940 28.540 56.340 ;
        RECT 28.840 54.940 30.540 56.340 ;
        RECT 30.840 54.940 32.540 56.340 ;
        RECT 32.840 54.940 34.540 56.340 ;
        RECT 34.840 54.940 36.540 56.340 ;
        RECT 36.840 54.940 38.540 56.340 ;
        RECT 38.840 54.940 40.540 56.340 ;
        RECT 40.840 54.940 42.540 56.340 ;
        RECT 42.840 54.940 44.540 56.340 ;
        RECT 44.840 54.940 46.540 56.340 ;
        RECT 46.840 54.940 48.540 56.340 ;
        RECT 48.840 54.940 50.540 56.340 ;
        RECT 50.840 54.940 52.540 56.340 ;
        RECT 52.840 54.940 54.540 56.340 ;
        RECT 54.840 54.940 56.540 56.340 ;
        RECT 56.840 54.940 58.540 56.340 ;
        RECT 58.840 54.940 60.540 56.340 ;
        RECT 60.840 54.940 62.540 56.340 ;
        RECT 62.840 54.940 64.540 56.340 ;
        RECT 64.840 54.940 66.540 56.340 ;
        RECT 66.840 54.940 68.540 56.340 ;
        RECT 68.840 54.940 70.540 56.340 ;
        RECT 70.840 54.940 72.540 56.340 ;
        RECT 72.840 54.940 74.540 56.340 ;
        RECT 86.575 54.940 88.275 56.340 ;
        RECT 88.575 54.940 90.275 56.340 ;
        RECT 90.575 54.940 92.275 56.340 ;
        RECT 92.575 54.940 94.275 56.340 ;
        RECT 94.575 54.940 96.275 56.340 ;
        RECT 96.575 54.940 98.275 56.340 ;
        RECT 98.575 54.940 100.275 56.340 ;
        RECT 100.575 54.940 102.275 56.340 ;
        RECT 102.575 54.940 104.275 56.340 ;
        RECT 104.575 54.940 106.275 56.340 ;
        RECT 106.575 54.940 108.275 56.340 ;
        RECT 108.575 54.940 110.275 56.340 ;
        RECT 110.575 54.940 112.275 56.340 ;
        RECT 112.575 54.940 114.275 56.340 ;
        RECT 114.575 54.940 116.275 56.340 ;
        RECT 116.575 54.940 118.275 56.340 ;
        RECT 118.575 54.940 120.275 56.340 ;
        RECT 120.575 54.940 122.275 56.340 ;
        RECT 122.575 54.940 124.275 56.340 ;
        RECT 124.575 54.940 126.275 56.340 ;
        RECT 126.575 54.940 128.275 56.340 ;
        RECT 128.575 54.940 130.275 56.340 ;
        RECT 130.575 54.940 132.275 56.340 ;
        RECT 132.575 54.940 134.275 56.340 ;
        RECT 134.575 54.940 136.275 56.340 ;
        RECT 136.575 54.940 138.275 56.340 ;
        RECT 138.575 54.940 140.275 56.340 ;
        RECT 140.575 54.940 142.275 56.340 ;
        RECT 142.575 54.940 144.275 56.340 ;
        RECT 144.575 54.940 146.275 56.340 ;
        RECT 146.575 54.940 148.275 56.340 ;
        RECT 148.575 54.940 150.275 56.340 ;
        RECT 150.575 54.940 152.275 56.340 ;
        RECT 152.575 54.940 154.275 56.340 ;
        RECT 6.840 53.090 8.540 54.490 ;
        RECT 8.840 53.090 10.540 54.490 ;
        RECT 10.840 53.090 12.540 54.490 ;
        RECT 12.840 53.090 14.540 54.490 ;
        RECT 14.840 53.090 16.540 54.490 ;
        RECT 16.840 53.090 18.540 54.490 ;
        RECT 18.840 53.090 20.540 54.490 ;
        RECT 20.840 53.090 22.540 54.490 ;
        RECT 22.840 53.090 24.540 54.490 ;
        RECT 24.840 53.090 26.540 54.490 ;
        RECT 26.840 53.090 28.540 54.490 ;
        RECT 28.840 53.090 30.540 54.490 ;
        RECT 30.840 53.090 32.540 54.490 ;
        RECT 32.840 53.090 34.540 54.490 ;
        RECT 34.840 53.090 36.540 54.490 ;
        RECT 36.840 53.090 38.540 54.490 ;
        RECT 38.840 53.090 40.540 54.490 ;
        RECT 40.840 53.090 42.540 54.490 ;
        RECT 42.840 53.090 44.540 54.490 ;
        RECT 44.840 53.090 46.540 54.490 ;
        RECT 46.840 53.090 48.540 54.490 ;
        RECT 48.840 53.090 50.540 54.490 ;
        RECT 50.840 53.090 52.540 54.490 ;
        RECT 52.840 53.090 54.540 54.490 ;
        RECT 54.840 53.090 56.540 54.490 ;
        RECT 56.840 53.090 58.540 54.490 ;
        RECT 58.840 53.090 60.540 54.490 ;
        RECT 60.840 53.090 62.540 54.490 ;
        RECT 62.840 53.090 64.540 54.490 ;
        RECT 64.840 53.090 66.540 54.490 ;
        RECT 66.840 53.090 68.540 54.490 ;
        RECT 68.840 53.090 70.540 54.490 ;
        RECT 70.840 53.090 72.540 54.490 ;
        RECT 72.840 53.090 74.540 54.490 ;
        RECT 86.575 53.090 88.275 54.490 ;
        RECT 88.575 53.090 90.275 54.490 ;
        RECT 90.575 53.090 92.275 54.490 ;
        RECT 92.575 53.090 94.275 54.490 ;
        RECT 94.575 53.090 96.275 54.490 ;
        RECT 96.575 53.090 98.275 54.490 ;
        RECT 98.575 53.090 100.275 54.490 ;
        RECT 100.575 53.090 102.275 54.490 ;
        RECT 102.575 53.090 104.275 54.490 ;
        RECT 104.575 53.090 106.275 54.490 ;
        RECT 106.575 53.090 108.275 54.490 ;
        RECT 108.575 53.090 110.275 54.490 ;
        RECT 110.575 53.090 112.275 54.490 ;
        RECT 112.575 53.090 114.275 54.490 ;
        RECT 114.575 53.090 116.275 54.490 ;
        RECT 116.575 53.090 118.275 54.490 ;
        RECT 118.575 53.090 120.275 54.490 ;
        RECT 120.575 53.090 122.275 54.490 ;
        RECT 122.575 53.090 124.275 54.490 ;
        RECT 124.575 53.090 126.275 54.490 ;
        RECT 126.575 53.090 128.275 54.490 ;
        RECT 128.575 53.090 130.275 54.490 ;
        RECT 130.575 53.090 132.275 54.490 ;
        RECT 132.575 53.090 134.275 54.490 ;
        RECT 134.575 53.090 136.275 54.490 ;
        RECT 136.575 53.090 138.275 54.490 ;
        RECT 138.575 53.090 140.275 54.490 ;
        RECT 140.575 53.090 142.275 54.490 ;
        RECT 142.575 53.090 144.275 54.490 ;
        RECT 144.575 53.090 146.275 54.490 ;
        RECT 146.575 53.090 148.275 54.490 ;
        RECT 148.575 53.090 150.275 54.490 ;
        RECT 150.575 53.090 152.275 54.490 ;
        RECT 152.575 53.090 154.275 54.490 ;
        RECT 6.840 51.240 8.540 52.640 ;
        RECT 8.840 51.240 10.540 52.640 ;
        RECT 10.840 51.240 12.540 52.640 ;
        RECT 12.840 51.240 14.540 52.640 ;
        RECT 14.840 51.240 16.540 52.640 ;
        RECT 16.840 51.240 18.540 52.640 ;
        RECT 18.840 51.240 20.540 52.640 ;
        RECT 20.840 51.240 22.540 52.640 ;
        RECT 22.840 51.240 24.540 52.640 ;
        RECT 24.840 51.240 26.540 52.640 ;
        RECT 26.840 51.240 28.540 52.640 ;
        RECT 28.840 51.240 30.540 52.640 ;
        RECT 30.840 51.240 32.540 52.640 ;
        RECT 32.840 51.240 34.540 52.640 ;
        RECT 34.840 51.240 36.540 52.640 ;
        RECT 36.840 51.240 38.540 52.640 ;
        RECT 38.840 51.240 40.540 52.640 ;
        RECT 40.840 51.240 42.540 52.640 ;
        RECT 42.840 51.240 44.540 52.640 ;
        RECT 44.840 51.240 46.540 52.640 ;
        RECT 46.840 51.240 48.540 52.640 ;
        RECT 48.840 51.240 50.540 52.640 ;
        RECT 50.840 51.240 52.540 52.640 ;
        RECT 52.840 51.240 54.540 52.640 ;
        RECT 54.840 51.240 56.540 52.640 ;
        RECT 56.840 51.240 58.540 52.640 ;
        RECT 58.840 51.240 60.540 52.640 ;
        RECT 60.840 51.240 62.540 52.640 ;
        RECT 62.840 51.240 64.540 52.640 ;
        RECT 64.840 51.240 66.540 52.640 ;
        RECT 66.840 51.240 68.540 52.640 ;
        RECT 68.840 51.240 70.540 52.640 ;
        RECT 70.840 51.240 72.540 52.640 ;
        RECT 72.840 51.240 74.540 52.640 ;
        RECT 86.575 51.240 88.275 52.640 ;
        RECT 88.575 51.240 90.275 52.640 ;
        RECT 90.575 51.240 92.275 52.640 ;
        RECT 92.575 51.240 94.275 52.640 ;
        RECT 94.575 51.240 96.275 52.640 ;
        RECT 96.575 51.240 98.275 52.640 ;
        RECT 98.575 51.240 100.275 52.640 ;
        RECT 100.575 51.240 102.275 52.640 ;
        RECT 102.575 51.240 104.275 52.640 ;
        RECT 104.575 51.240 106.275 52.640 ;
        RECT 106.575 51.240 108.275 52.640 ;
        RECT 108.575 51.240 110.275 52.640 ;
        RECT 110.575 51.240 112.275 52.640 ;
        RECT 112.575 51.240 114.275 52.640 ;
        RECT 114.575 51.240 116.275 52.640 ;
        RECT 116.575 51.240 118.275 52.640 ;
        RECT 118.575 51.240 120.275 52.640 ;
        RECT 120.575 51.240 122.275 52.640 ;
        RECT 122.575 51.240 124.275 52.640 ;
        RECT 124.575 51.240 126.275 52.640 ;
        RECT 126.575 51.240 128.275 52.640 ;
        RECT 128.575 51.240 130.275 52.640 ;
        RECT 130.575 51.240 132.275 52.640 ;
        RECT 132.575 51.240 134.275 52.640 ;
        RECT 134.575 51.240 136.275 52.640 ;
        RECT 136.575 51.240 138.275 52.640 ;
        RECT 138.575 51.240 140.275 52.640 ;
        RECT 140.575 51.240 142.275 52.640 ;
        RECT 142.575 51.240 144.275 52.640 ;
        RECT 144.575 51.240 146.275 52.640 ;
        RECT 146.575 51.240 148.275 52.640 ;
        RECT 148.575 51.240 150.275 52.640 ;
        RECT 150.575 51.240 152.275 52.640 ;
        RECT 152.575 51.240 154.275 52.640 ;
        RECT 6.840 49.390 8.540 50.790 ;
        RECT 8.840 49.390 10.540 50.790 ;
        RECT 10.840 49.390 12.540 50.790 ;
        RECT 12.840 49.390 14.540 50.790 ;
        RECT 14.840 49.390 16.540 50.790 ;
        RECT 16.840 49.390 18.540 50.790 ;
        RECT 18.840 49.390 20.540 50.790 ;
        RECT 20.840 49.390 22.540 50.790 ;
        RECT 22.840 49.390 24.540 50.790 ;
        RECT 24.840 49.390 26.540 50.790 ;
        RECT 26.840 49.390 28.540 50.790 ;
        RECT 28.840 49.390 30.540 50.790 ;
        RECT 30.840 49.390 32.540 50.790 ;
        RECT 32.840 49.390 34.540 50.790 ;
        RECT 34.840 49.390 36.540 50.790 ;
        RECT 36.840 49.390 38.540 50.790 ;
        RECT 38.840 49.390 40.540 50.790 ;
        RECT 40.840 49.390 42.540 50.790 ;
        RECT 42.840 49.390 44.540 50.790 ;
        RECT 44.840 49.390 46.540 50.790 ;
        RECT 46.840 49.390 48.540 50.790 ;
        RECT 48.840 49.390 50.540 50.790 ;
        RECT 50.840 49.390 52.540 50.790 ;
        RECT 52.840 49.390 54.540 50.790 ;
        RECT 54.840 49.390 56.540 50.790 ;
        RECT 56.840 49.390 58.540 50.790 ;
        RECT 58.840 49.390 60.540 50.790 ;
        RECT 60.840 49.390 62.540 50.790 ;
        RECT 62.840 49.390 64.540 50.790 ;
        RECT 64.840 49.390 66.540 50.790 ;
        RECT 66.840 49.390 68.540 50.790 ;
        RECT 68.840 49.390 70.540 50.790 ;
        RECT 70.840 49.390 72.540 50.790 ;
        RECT 72.840 49.390 74.540 50.790 ;
        RECT 86.575 49.390 88.275 50.790 ;
        RECT 88.575 49.390 90.275 50.790 ;
        RECT 90.575 49.390 92.275 50.790 ;
        RECT 92.575 49.390 94.275 50.790 ;
        RECT 94.575 49.390 96.275 50.790 ;
        RECT 96.575 49.390 98.275 50.790 ;
        RECT 98.575 49.390 100.275 50.790 ;
        RECT 100.575 49.390 102.275 50.790 ;
        RECT 102.575 49.390 104.275 50.790 ;
        RECT 104.575 49.390 106.275 50.790 ;
        RECT 106.575 49.390 108.275 50.790 ;
        RECT 108.575 49.390 110.275 50.790 ;
        RECT 110.575 49.390 112.275 50.790 ;
        RECT 112.575 49.390 114.275 50.790 ;
        RECT 114.575 49.390 116.275 50.790 ;
        RECT 116.575 49.390 118.275 50.790 ;
        RECT 118.575 49.390 120.275 50.790 ;
        RECT 120.575 49.390 122.275 50.790 ;
        RECT 122.575 49.390 124.275 50.790 ;
        RECT 124.575 49.390 126.275 50.790 ;
        RECT 126.575 49.390 128.275 50.790 ;
        RECT 128.575 49.390 130.275 50.790 ;
        RECT 130.575 49.390 132.275 50.790 ;
        RECT 132.575 49.390 134.275 50.790 ;
        RECT 134.575 49.390 136.275 50.790 ;
        RECT 136.575 49.390 138.275 50.790 ;
        RECT 138.575 49.390 140.275 50.790 ;
        RECT 140.575 49.390 142.275 50.790 ;
        RECT 142.575 49.390 144.275 50.790 ;
        RECT 144.575 49.390 146.275 50.790 ;
        RECT 146.575 49.390 148.275 50.790 ;
        RECT 148.575 49.390 150.275 50.790 ;
        RECT 150.575 49.390 152.275 50.790 ;
        RECT 152.575 49.390 154.275 50.790 ;
        RECT 6.840 47.540 8.540 48.940 ;
        RECT 8.840 47.540 10.540 48.940 ;
        RECT 10.840 47.540 12.540 48.940 ;
        RECT 12.840 47.540 14.540 48.940 ;
        RECT 14.840 47.540 16.540 48.940 ;
        RECT 16.840 47.540 18.540 48.940 ;
        RECT 18.840 47.540 20.540 48.940 ;
        RECT 20.840 47.540 22.540 48.940 ;
        RECT 22.840 47.540 24.540 48.940 ;
        RECT 24.840 47.540 26.540 48.940 ;
        RECT 26.840 47.540 28.540 48.940 ;
        RECT 28.840 47.540 30.540 48.940 ;
        RECT 30.840 47.540 32.540 48.940 ;
        RECT 32.840 47.540 34.540 48.940 ;
        RECT 34.840 47.540 36.540 48.940 ;
        RECT 36.840 47.540 38.540 48.940 ;
        RECT 38.840 47.540 40.540 48.940 ;
        RECT 40.840 47.540 42.540 48.940 ;
        RECT 42.840 47.540 44.540 48.940 ;
        RECT 44.840 47.540 46.540 48.940 ;
        RECT 46.840 47.540 48.540 48.940 ;
        RECT 48.840 47.540 50.540 48.940 ;
        RECT 50.840 47.540 52.540 48.940 ;
        RECT 52.840 47.540 54.540 48.940 ;
        RECT 54.840 47.540 56.540 48.940 ;
        RECT 56.840 47.540 58.540 48.940 ;
        RECT 58.840 47.540 60.540 48.940 ;
        RECT 60.840 47.540 62.540 48.940 ;
        RECT 62.840 47.540 64.540 48.940 ;
        RECT 64.840 47.540 66.540 48.940 ;
        RECT 66.840 47.540 68.540 48.940 ;
        RECT 68.840 47.540 70.540 48.940 ;
        RECT 70.840 47.540 72.540 48.940 ;
        RECT 72.840 47.540 74.540 48.940 ;
        RECT 86.575 47.540 88.275 48.940 ;
        RECT 88.575 47.540 90.275 48.940 ;
        RECT 90.575 47.540 92.275 48.940 ;
        RECT 92.575 47.540 94.275 48.940 ;
        RECT 94.575 47.540 96.275 48.940 ;
        RECT 96.575 47.540 98.275 48.940 ;
        RECT 98.575 47.540 100.275 48.940 ;
        RECT 100.575 47.540 102.275 48.940 ;
        RECT 102.575 47.540 104.275 48.940 ;
        RECT 104.575 47.540 106.275 48.940 ;
        RECT 106.575 47.540 108.275 48.940 ;
        RECT 108.575 47.540 110.275 48.940 ;
        RECT 110.575 47.540 112.275 48.940 ;
        RECT 112.575 47.540 114.275 48.940 ;
        RECT 114.575 47.540 116.275 48.940 ;
        RECT 116.575 47.540 118.275 48.940 ;
        RECT 118.575 47.540 120.275 48.940 ;
        RECT 120.575 47.540 122.275 48.940 ;
        RECT 122.575 47.540 124.275 48.940 ;
        RECT 124.575 47.540 126.275 48.940 ;
        RECT 126.575 47.540 128.275 48.940 ;
        RECT 128.575 47.540 130.275 48.940 ;
        RECT 130.575 47.540 132.275 48.940 ;
        RECT 132.575 47.540 134.275 48.940 ;
        RECT 134.575 47.540 136.275 48.940 ;
        RECT 136.575 47.540 138.275 48.940 ;
        RECT 138.575 47.540 140.275 48.940 ;
        RECT 140.575 47.540 142.275 48.940 ;
        RECT 142.575 47.540 144.275 48.940 ;
        RECT 144.575 47.540 146.275 48.940 ;
        RECT 146.575 47.540 148.275 48.940 ;
        RECT 148.575 47.540 150.275 48.940 ;
        RECT 150.575 47.540 152.275 48.940 ;
        RECT 152.575 47.540 154.275 48.940 ;
        RECT 6.840 45.690 8.540 47.090 ;
        RECT 8.840 45.690 10.540 47.090 ;
        RECT 10.840 45.690 12.540 47.090 ;
        RECT 12.840 45.690 14.540 47.090 ;
        RECT 14.840 45.690 16.540 47.090 ;
        RECT 16.840 45.690 18.540 47.090 ;
        RECT 18.840 45.690 20.540 47.090 ;
        RECT 20.840 45.690 22.540 47.090 ;
        RECT 22.840 45.690 24.540 47.090 ;
        RECT 24.840 45.690 26.540 47.090 ;
        RECT 26.840 45.690 28.540 47.090 ;
        RECT 28.840 45.690 30.540 47.090 ;
        RECT 30.840 45.690 32.540 47.090 ;
        RECT 32.840 45.690 34.540 47.090 ;
        RECT 34.840 45.690 36.540 47.090 ;
        RECT 36.840 45.690 38.540 47.090 ;
        RECT 38.840 45.690 40.540 47.090 ;
        RECT 40.840 45.690 42.540 47.090 ;
        RECT 42.840 45.690 44.540 47.090 ;
        RECT 44.840 45.690 46.540 47.090 ;
        RECT 46.840 45.690 48.540 47.090 ;
        RECT 48.840 45.690 50.540 47.090 ;
        RECT 50.840 45.690 52.540 47.090 ;
        RECT 52.840 45.690 54.540 47.090 ;
        RECT 54.840 45.690 56.540 47.090 ;
        RECT 56.840 45.690 58.540 47.090 ;
        RECT 58.840 45.690 60.540 47.090 ;
        RECT 60.840 45.690 62.540 47.090 ;
        RECT 62.840 45.690 64.540 47.090 ;
        RECT 64.840 45.690 66.540 47.090 ;
        RECT 66.840 45.690 68.540 47.090 ;
        RECT 68.840 45.690 70.540 47.090 ;
        RECT 70.840 45.690 72.540 47.090 ;
        RECT 72.840 45.690 74.540 47.090 ;
        RECT 86.575 45.690 88.275 47.090 ;
        RECT 88.575 45.690 90.275 47.090 ;
        RECT 90.575 45.690 92.275 47.090 ;
        RECT 92.575 45.690 94.275 47.090 ;
        RECT 94.575 45.690 96.275 47.090 ;
        RECT 96.575 45.690 98.275 47.090 ;
        RECT 98.575 45.690 100.275 47.090 ;
        RECT 100.575 45.690 102.275 47.090 ;
        RECT 102.575 45.690 104.275 47.090 ;
        RECT 104.575 45.690 106.275 47.090 ;
        RECT 106.575 45.690 108.275 47.090 ;
        RECT 108.575 45.690 110.275 47.090 ;
        RECT 110.575 45.690 112.275 47.090 ;
        RECT 112.575 45.690 114.275 47.090 ;
        RECT 114.575 45.690 116.275 47.090 ;
        RECT 116.575 45.690 118.275 47.090 ;
        RECT 118.575 45.690 120.275 47.090 ;
        RECT 120.575 45.690 122.275 47.090 ;
        RECT 122.575 45.690 124.275 47.090 ;
        RECT 124.575 45.690 126.275 47.090 ;
        RECT 126.575 45.690 128.275 47.090 ;
        RECT 128.575 45.690 130.275 47.090 ;
        RECT 130.575 45.690 132.275 47.090 ;
        RECT 132.575 45.690 134.275 47.090 ;
        RECT 134.575 45.690 136.275 47.090 ;
        RECT 136.575 45.690 138.275 47.090 ;
        RECT 138.575 45.690 140.275 47.090 ;
        RECT 140.575 45.690 142.275 47.090 ;
        RECT 142.575 45.690 144.275 47.090 ;
        RECT 144.575 45.690 146.275 47.090 ;
        RECT 146.575 45.690 148.275 47.090 ;
        RECT 148.575 45.690 150.275 47.090 ;
        RECT 150.575 45.690 152.275 47.090 ;
        RECT 152.575 45.690 154.275 47.090 ;
        RECT 6.840 43.840 8.540 45.240 ;
        RECT 8.840 43.840 10.540 45.240 ;
        RECT 10.840 43.840 12.540 45.240 ;
        RECT 12.840 43.840 14.540 45.240 ;
        RECT 14.840 43.840 16.540 45.240 ;
        RECT 16.840 43.840 18.540 45.240 ;
        RECT 18.840 43.840 20.540 45.240 ;
        RECT 20.840 43.840 22.540 45.240 ;
        RECT 22.840 43.840 24.540 45.240 ;
        RECT 24.840 43.840 26.540 45.240 ;
        RECT 26.840 43.840 28.540 45.240 ;
        RECT 28.840 43.840 30.540 45.240 ;
        RECT 30.840 43.840 32.540 45.240 ;
        RECT 32.840 43.840 34.540 45.240 ;
        RECT 34.840 43.840 36.540 45.240 ;
        RECT 36.840 43.840 38.540 45.240 ;
        RECT 38.840 43.840 40.540 45.240 ;
        RECT 40.840 43.840 42.540 45.240 ;
        RECT 42.840 43.840 44.540 45.240 ;
        RECT 44.840 43.840 46.540 45.240 ;
        RECT 46.840 43.840 48.540 45.240 ;
        RECT 48.840 43.840 50.540 45.240 ;
        RECT 50.840 43.840 52.540 45.240 ;
        RECT 52.840 43.840 54.540 45.240 ;
        RECT 54.840 43.840 56.540 45.240 ;
        RECT 56.840 43.840 58.540 45.240 ;
        RECT 58.840 43.840 60.540 45.240 ;
        RECT 60.840 43.840 62.540 45.240 ;
        RECT 62.840 43.840 64.540 45.240 ;
        RECT 64.840 43.840 66.540 45.240 ;
        RECT 66.840 43.840 68.540 45.240 ;
        RECT 68.840 43.840 70.540 45.240 ;
        RECT 70.840 43.840 72.540 45.240 ;
        RECT 72.840 43.840 74.540 45.240 ;
        RECT 86.575 43.840 88.275 45.240 ;
        RECT 88.575 43.840 90.275 45.240 ;
        RECT 90.575 43.840 92.275 45.240 ;
        RECT 92.575 43.840 94.275 45.240 ;
        RECT 94.575 43.840 96.275 45.240 ;
        RECT 96.575 43.840 98.275 45.240 ;
        RECT 98.575 43.840 100.275 45.240 ;
        RECT 100.575 43.840 102.275 45.240 ;
        RECT 102.575 43.840 104.275 45.240 ;
        RECT 104.575 43.840 106.275 45.240 ;
        RECT 106.575 43.840 108.275 45.240 ;
        RECT 108.575 43.840 110.275 45.240 ;
        RECT 110.575 43.840 112.275 45.240 ;
        RECT 112.575 43.840 114.275 45.240 ;
        RECT 114.575 43.840 116.275 45.240 ;
        RECT 116.575 43.840 118.275 45.240 ;
        RECT 118.575 43.840 120.275 45.240 ;
        RECT 120.575 43.840 122.275 45.240 ;
        RECT 122.575 43.840 124.275 45.240 ;
        RECT 124.575 43.840 126.275 45.240 ;
        RECT 126.575 43.840 128.275 45.240 ;
        RECT 128.575 43.840 130.275 45.240 ;
        RECT 130.575 43.840 132.275 45.240 ;
        RECT 132.575 43.840 134.275 45.240 ;
        RECT 134.575 43.840 136.275 45.240 ;
        RECT 136.575 43.840 138.275 45.240 ;
        RECT 138.575 43.840 140.275 45.240 ;
        RECT 140.575 43.840 142.275 45.240 ;
        RECT 142.575 43.840 144.275 45.240 ;
        RECT 144.575 43.840 146.275 45.240 ;
        RECT 146.575 43.840 148.275 45.240 ;
        RECT 148.575 43.840 150.275 45.240 ;
        RECT 150.575 43.840 152.275 45.240 ;
        RECT 152.575 43.840 154.275 45.240 ;
        RECT 6.840 41.990 8.540 43.390 ;
        RECT 8.840 41.990 10.540 43.390 ;
        RECT 10.840 41.990 12.540 43.390 ;
        RECT 12.840 41.990 14.540 43.390 ;
        RECT 14.840 41.990 16.540 43.390 ;
        RECT 16.840 41.990 18.540 43.390 ;
        RECT 18.840 41.990 20.540 43.390 ;
        RECT 20.840 41.990 22.540 43.390 ;
        RECT 22.840 41.990 24.540 43.390 ;
        RECT 24.840 41.990 26.540 43.390 ;
        RECT 26.840 41.990 28.540 43.390 ;
        RECT 28.840 41.990 30.540 43.390 ;
        RECT 30.840 41.990 32.540 43.390 ;
        RECT 32.840 41.990 34.540 43.390 ;
        RECT 34.840 41.990 36.540 43.390 ;
        RECT 36.840 41.990 38.540 43.390 ;
        RECT 38.840 41.990 40.540 43.390 ;
        RECT 40.840 41.990 42.540 43.390 ;
        RECT 42.840 41.990 44.540 43.390 ;
        RECT 44.840 41.990 46.540 43.390 ;
        RECT 46.840 41.990 48.540 43.390 ;
        RECT 48.840 41.990 50.540 43.390 ;
        RECT 50.840 41.990 52.540 43.390 ;
        RECT 52.840 41.990 54.540 43.390 ;
        RECT 54.840 41.990 56.540 43.390 ;
        RECT 56.840 41.990 58.540 43.390 ;
        RECT 58.840 41.990 60.540 43.390 ;
        RECT 60.840 41.990 62.540 43.390 ;
        RECT 62.840 41.990 64.540 43.390 ;
        RECT 64.840 41.990 66.540 43.390 ;
        RECT 66.840 41.990 68.540 43.390 ;
        RECT 68.840 41.990 70.540 43.390 ;
        RECT 70.840 41.990 72.540 43.390 ;
        RECT 72.840 41.990 74.540 43.390 ;
        RECT 86.575 41.990 88.275 43.390 ;
        RECT 88.575 41.990 90.275 43.390 ;
        RECT 90.575 41.990 92.275 43.390 ;
        RECT 92.575 41.990 94.275 43.390 ;
        RECT 94.575 41.990 96.275 43.390 ;
        RECT 96.575 41.990 98.275 43.390 ;
        RECT 98.575 41.990 100.275 43.390 ;
        RECT 100.575 41.990 102.275 43.390 ;
        RECT 102.575 41.990 104.275 43.390 ;
        RECT 104.575 41.990 106.275 43.390 ;
        RECT 106.575 41.990 108.275 43.390 ;
        RECT 108.575 41.990 110.275 43.390 ;
        RECT 110.575 41.990 112.275 43.390 ;
        RECT 112.575 41.990 114.275 43.390 ;
        RECT 114.575 41.990 116.275 43.390 ;
        RECT 116.575 41.990 118.275 43.390 ;
        RECT 118.575 41.990 120.275 43.390 ;
        RECT 120.575 41.990 122.275 43.390 ;
        RECT 122.575 41.990 124.275 43.390 ;
        RECT 124.575 41.990 126.275 43.390 ;
        RECT 126.575 41.990 128.275 43.390 ;
        RECT 128.575 41.990 130.275 43.390 ;
        RECT 130.575 41.990 132.275 43.390 ;
        RECT 132.575 41.990 134.275 43.390 ;
        RECT 134.575 41.990 136.275 43.390 ;
        RECT 136.575 41.990 138.275 43.390 ;
        RECT 138.575 41.990 140.275 43.390 ;
        RECT 140.575 41.990 142.275 43.390 ;
        RECT 142.575 41.990 144.275 43.390 ;
        RECT 144.575 41.990 146.275 43.390 ;
        RECT 146.575 41.990 148.275 43.390 ;
        RECT 148.575 41.990 150.275 43.390 ;
        RECT 150.575 41.990 152.275 43.390 ;
        RECT 152.575 41.990 154.275 43.390 ;
        RECT 6.840 40.140 8.540 41.540 ;
        RECT 8.840 40.140 10.540 41.540 ;
        RECT 10.840 40.140 12.540 41.540 ;
        RECT 12.840 40.140 14.540 41.540 ;
        RECT 14.840 40.140 16.540 41.540 ;
        RECT 16.840 40.140 18.540 41.540 ;
        RECT 18.840 40.140 20.540 41.540 ;
        RECT 20.840 40.140 22.540 41.540 ;
        RECT 22.840 40.140 24.540 41.540 ;
        RECT 24.840 40.140 26.540 41.540 ;
        RECT 26.840 40.140 28.540 41.540 ;
        RECT 28.840 40.140 30.540 41.540 ;
        RECT 30.840 40.140 32.540 41.540 ;
        RECT 32.840 40.140 34.540 41.540 ;
        RECT 34.840 40.140 36.540 41.540 ;
        RECT 36.840 40.140 38.540 41.540 ;
        RECT 38.840 40.140 40.540 41.540 ;
        RECT 40.840 40.140 42.540 41.540 ;
        RECT 42.840 40.140 44.540 41.540 ;
        RECT 44.840 40.140 46.540 41.540 ;
        RECT 46.840 40.140 48.540 41.540 ;
        RECT 48.840 40.140 50.540 41.540 ;
        RECT 50.840 40.140 52.540 41.540 ;
        RECT 52.840 40.140 54.540 41.540 ;
        RECT 54.840 40.140 56.540 41.540 ;
        RECT 56.840 40.140 58.540 41.540 ;
        RECT 58.840 40.140 60.540 41.540 ;
        RECT 60.840 40.140 62.540 41.540 ;
        RECT 62.840 40.140 64.540 41.540 ;
        RECT 64.840 40.140 66.540 41.540 ;
        RECT 66.840 40.140 68.540 41.540 ;
        RECT 68.840 40.140 70.540 41.540 ;
        RECT 70.840 40.140 72.540 41.540 ;
        RECT 72.840 40.140 74.540 41.540 ;
        RECT 86.575 40.140 88.275 41.540 ;
        RECT 88.575 40.140 90.275 41.540 ;
        RECT 90.575 40.140 92.275 41.540 ;
        RECT 92.575 40.140 94.275 41.540 ;
        RECT 94.575 40.140 96.275 41.540 ;
        RECT 96.575 40.140 98.275 41.540 ;
        RECT 98.575 40.140 100.275 41.540 ;
        RECT 100.575 40.140 102.275 41.540 ;
        RECT 102.575 40.140 104.275 41.540 ;
        RECT 104.575 40.140 106.275 41.540 ;
        RECT 106.575 40.140 108.275 41.540 ;
        RECT 108.575 40.140 110.275 41.540 ;
        RECT 110.575 40.140 112.275 41.540 ;
        RECT 112.575 40.140 114.275 41.540 ;
        RECT 114.575 40.140 116.275 41.540 ;
        RECT 116.575 40.140 118.275 41.540 ;
        RECT 118.575 40.140 120.275 41.540 ;
        RECT 120.575 40.140 122.275 41.540 ;
        RECT 122.575 40.140 124.275 41.540 ;
        RECT 124.575 40.140 126.275 41.540 ;
        RECT 126.575 40.140 128.275 41.540 ;
        RECT 128.575 40.140 130.275 41.540 ;
        RECT 130.575 40.140 132.275 41.540 ;
        RECT 132.575 40.140 134.275 41.540 ;
        RECT 134.575 40.140 136.275 41.540 ;
        RECT 136.575 40.140 138.275 41.540 ;
        RECT 138.575 40.140 140.275 41.540 ;
        RECT 140.575 40.140 142.275 41.540 ;
        RECT 142.575 40.140 144.275 41.540 ;
        RECT 144.575 40.140 146.275 41.540 ;
        RECT 146.575 40.140 148.275 41.540 ;
        RECT 148.575 40.140 150.275 41.540 ;
        RECT 150.575 40.140 152.275 41.540 ;
        RECT 152.575 40.140 154.275 41.540 ;
        RECT 6.840 38.290 8.540 39.690 ;
        RECT 8.840 38.290 10.540 39.690 ;
        RECT 10.840 38.290 12.540 39.690 ;
        RECT 12.840 38.290 14.540 39.690 ;
        RECT 14.840 38.290 16.540 39.690 ;
        RECT 16.840 38.290 18.540 39.690 ;
        RECT 18.840 38.290 20.540 39.690 ;
        RECT 20.840 38.290 22.540 39.690 ;
        RECT 22.840 38.290 24.540 39.690 ;
        RECT 24.840 38.290 26.540 39.690 ;
        RECT 26.840 38.290 28.540 39.690 ;
        RECT 28.840 38.290 30.540 39.690 ;
        RECT 30.840 38.290 32.540 39.690 ;
        RECT 32.840 38.290 34.540 39.690 ;
        RECT 34.840 38.290 36.540 39.690 ;
        RECT 36.840 38.290 38.540 39.690 ;
        RECT 38.840 38.290 40.540 39.690 ;
        RECT 40.840 38.290 42.540 39.690 ;
        RECT 42.840 38.290 44.540 39.690 ;
        RECT 44.840 38.290 46.540 39.690 ;
        RECT 46.840 38.290 48.540 39.690 ;
        RECT 48.840 38.290 50.540 39.690 ;
        RECT 50.840 38.290 52.540 39.690 ;
        RECT 52.840 38.290 54.540 39.690 ;
        RECT 54.840 38.290 56.540 39.690 ;
        RECT 56.840 38.290 58.540 39.690 ;
        RECT 58.840 38.290 60.540 39.690 ;
        RECT 60.840 38.290 62.540 39.690 ;
        RECT 62.840 38.290 64.540 39.690 ;
        RECT 64.840 38.290 66.540 39.690 ;
        RECT 66.840 38.290 68.540 39.690 ;
        RECT 68.840 38.290 70.540 39.690 ;
        RECT 70.840 38.290 72.540 39.690 ;
        RECT 72.840 38.290 74.540 39.690 ;
        RECT 86.575 38.290 88.275 39.690 ;
        RECT 88.575 38.290 90.275 39.690 ;
        RECT 90.575 38.290 92.275 39.690 ;
        RECT 92.575 38.290 94.275 39.690 ;
        RECT 94.575 38.290 96.275 39.690 ;
        RECT 96.575 38.290 98.275 39.690 ;
        RECT 98.575 38.290 100.275 39.690 ;
        RECT 100.575 38.290 102.275 39.690 ;
        RECT 102.575 38.290 104.275 39.690 ;
        RECT 104.575 38.290 106.275 39.690 ;
        RECT 106.575 38.290 108.275 39.690 ;
        RECT 108.575 38.290 110.275 39.690 ;
        RECT 110.575 38.290 112.275 39.690 ;
        RECT 112.575 38.290 114.275 39.690 ;
        RECT 114.575 38.290 116.275 39.690 ;
        RECT 116.575 38.290 118.275 39.690 ;
        RECT 118.575 38.290 120.275 39.690 ;
        RECT 120.575 38.290 122.275 39.690 ;
        RECT 122.575 38.290 124.275 39.690 ;
        RECT 124.575 38.290 126.275 39.690 ;
        RECT 126.575 38.290 128.275 39.690 ;
        RECT 128.575 38.290 130.275 39.690 ;
        RECT 130.575 38.290 132.275 39.690 ;
        RECT 132.575 38.290 134.275 39.690 ;
        RECT 134.575 38.290 136.275 39.690 ;
        RECT 136.575 38.290 138.275 39.690 ;
        RECT 138.575 38.290 140.275 39.690 ;
        RECT 140.575 38.290 142.275 39.690 ;
        RECT 142.575 38.290 144.275 39.690 ;
        RECT 144.575 38.290 146.275 39.690 ;
        RECT 146.575 38.290 148.275 39.690 ;
        RECT 148.575 38.290 150.275 39.690 ;
        RECT 150.575 38.290 152.275 39.690 ;
        RECT 152.575 38.290 154.275 39.690 ;
        RECT 6.840 36.440 8.540 37.840 ;
        RECT 8.840 36.440 10.540 37.840 ;
        RECT 10.840 36.440 12.540 37.840 ;
        RECT 12.840 36.440 14.540 37.840 ;
        RECT 14.840 36.440 16.540 37.840 ;
        RECT 16.840 36.440 18.540 37.840 ;
        RECT 18.840 36.440 20.540 37.840 ;
        RECT 20.840 36.440 22.540 37.840 ;
        RECT 22.840 36.440 24.540 37.840 ;
        RECT 24.840 36.440 26.540 37.840 ;
        RECT 26.840 36.440 28.540 37.840 ;
        RECT 28.840 36.440 30.540 37.840 ;
        RECT 30.840 36.440 32.540 37.840 ;
        RECT 32.840 36.440 34.540 37.840 ;
        RECT 34.840 36.440 36.540 37.840 ;
        RECT 36.840 36.440 38.540 37.840 ;
        RECT 38.840 36.440 40.540 37.840 ;
        RECT 40.840 36.440 42.540 37.840 ;
        RECT 42.840 36.440 44.540 37.840 ;
        RECT 44.840 36.440 46.540 37.840 ;
        RECT 46.840 36.440 48.540 37.840 ;
        RECT 48.840 36.440 50.540 37.840 ;
        RECT 50.840 36.440 52.540 37.840 ;
        RECT 52.840 36.440 54.540 37.840 ;
        RECT 54.840 36.440 56.540 37.840 ;
        RECT 56.840 36.440 58.540 37.840 ;
        RECT 58.840 36.440 60.540 37.840 ;
        RECT 60.840 36.440 62.540 37.840 ;
        RECT 62.840 36.440 64.540 37.840 ;
        RECT 64.840 36.440 66.540 37.840 ;
        RECT 66.840 36.440 68.540 37.840 ;
        RECT 68.840 36.440 70.540 37.840 ;
        RECT 70.840 36.440 72.540 37.840 ;
        RECT 72.840 36.440 74.540 37.840 ;
        RECT 86.575 36.440 88.275 37.840 ;
        RECT 88.575 36.440 90.275 37.840 ;
        RECT 90.575 36.440 92.275 37.840 ;
        RECT 92.575 36.440 94.275 37.840 ;
        RECT 94.575 36.440 96.275 37.840 ;
        RECT 96.575 36.440 98.275 37.840 ;
        RECT 98.575 36.440 100.275 37.840 ;
        RECT 100.575 36.440 102.275 37.840 ;
        RECT 102.575 36.440 104.275 37.840 ;
        RECT 104.575 36.440 106.275 37.840 ;
        RECT 106.575 36.440 108.275 37.840 ;
        RECT 108.575 36.440 110.275 37.840 ;
        RECT 110.575 36.440 112.275 37.840 ;
        RECT 112.575 36.440 114.275 37.840 ;
        RECT 114.575 36.440 116.275 37.840 ;
        RECT 116.575 36.440 118.275 37.840 ;
        RECT 118.575 36.440 120.275 37.840 ;
        RECT 120.575 36.440 122.275 37.840 ;
        RECT 122.575 36.440 124.275 37.840 ;
        RECT 124.575 36.440 126.275 37.840 ;
        RECT 126.575 36.440 128.275 37.840 ;
        RECT 128.575 36.440 130.275 37.840 ;
        RECT 130.575 36.440 132.275 37.840 ;
        RECT 132.575 36.440 134.275 37.840 ;
        RECT 134.575 36.440 136.275 37.840 ;
        RECT 136.575 36.440 138.275 37.840 ;
        RECT 138.575 36.440 140.275 37.840 ;
        RECT 140.575 36.440 142.275 37.840 ;
        RECT 142.575 36.440 144.275 37.840 ;
        RECT 144.575 36.440 146.275 37.840 ;
        RECT 146.575 36.440 148.275 37.840 ;
        RECT 148.575 36.440 150.275 37.840 ;
        RECT 150.575 36.440 152.275 37.840 ;
        RECT 152.575 36.440 154.275 37.840 ;
        RECT 6.840 34.590 8.540 35.990 ;
        RECT 8.840 34.590 10.540 35.990 ;
        RECT 10.840 34.590 12.540 35.990 ;
        RECT 12.840 34.590 14.540 35.990 ;
        RECT 14.840 34.590 16.540 35.990 ;
        RECT 16.840 34.590 18.540 35.990 ;
        RECT 18.840 34.590 20.540 35.990 ;
        RECT 20.840 34.590 22.540 35.990 ;
        RECT 22.840 34.590 24.540 35.990 ;
        RECT 24.840 34.590 26.540 35.990 ;
        RECT 26.840 34.590 28.540 35.990 ;
        RECT 28.840 34.590 30.540 35.990 ;
        RECT 30.840 34.590 32.540 35.990 ;
        RECT 32.840 34.590 34.540 35.990 ;
        RECT 34.840 34.590 36.540 35.990 ;
        RECT 36.840 34.590 38.540 35.990 ;
        RECT 38.840 34.590 40.540 35.990 ;
        RECT 40.840 34.590 42.540 35.990 ;
        RECT 42.840 34.590 44.540 35.990 ;
        RECT 44.840 34.590 46.540 35.990 ;
        RECT 46.840 34.590 48.540 35.990 ;
        RECT 48.840 34.590 50.540 35.990 ;
        RECT 50.840 34.590 52.540 35.990 ;
        RECT 52.840 34.590 54.540 35.990 ;
        RECT 54.840 34.590 56.540 35.990 ;
        RECT 56.840 34.590 58.540 35.990 ;
        RECT 58.840 34.590 60.540 35.990 ;
        RECT 60.840 34.590 62.540 35.990 ;
        RECT 62.840 34.590 64.540 35.990 ;
        RECT 64.840 34.590 66.540 35.990 ;
        RECT 66.840 34.590 68.540 35.990 ;
        RECT 68.840 34.590 70.540 35.990 ;
        RECT 70.840 34.590 72.540 35.990 ;
        RECT 72.840 34.590 74.540 35.990 ;
        RECT 86.575 34.590 88.275 35.990 ;
        RECT 88.575 34.590 90.275 35.990 ;
        RECT 90.575 34.590 92.275 35.990 ;
        RECT 92.575 34.590 94.275 35.990 ;
        RECT 94.575 34.590 96.275 35.990 ;
        RECT 96.575 34.590 98.275 35.990 ;
        RECT 98.575 34.590 100.275 35.990 ;
        RECT 100.575 34.590 102.275 35.990 ;
        RECT 102.575 34.590 104.275 35.990 ;
        RECT 104.575 34.590 106.275 35.990 ;
        RECT 106.575 34.590 108.275 35.990 ;
        RECT 108.575 34.590 110.275 35.990 ;
        RECT 110.575 34.590 112.275 35.990 ;
        RECT 112.575 34.590 114.275 35.990 ;
        RECT 114.575 34.590 116.275 35.990 ;
        RECT 116.575 34.590 118.275 35.990 ;
        RECT 118.575 34.590 120.275 35.990 ;
        RECT 120.575 34.590 122.275 35.990 ;
        RECT 122.575 34.590 124.275 35.990 ;
        RECT 124.575 34.590 126.275 35.990 ;
        RECT 126.575 34.590 128.275 35.990 ;
        RECT 128.575 34.590 130.275 35.990 ;
        RECT 130.575 34.590 132.275 35.990 ;
        RECT 132.575 34.590 134.275 35.990 ;
        RECT 134.575 34.590 136.275 35.990 ;
        RECT 136.575 34.590 138.275 35.990 ;
        RECT 138.575 34.590 140.275 35.990 ;
        RECT 140.575 34.590 142.275 35.990 ;
        RECT 142.575 34.590 144.275 35.990 ;
        RECT 144.575 34.590 146.275 35.990 ;
        RECT 146.575 34.590 148.275 35.990 ;
        RECT 148.575 34.590 150.275 35.990 ;
        RECT 150.575 34.590 152.275 35.990 ;
        RECT 152.575 34.590 154.275 35.990 ;
        RECT 6.840 32.740 8.540 34.140 ;
        RECT 8.840 32.740 10.540 34.140 ;
        RECT 10.840 32.740 12.540 34.140 ;
        RECT 12.840 32.740 14.540 34.140 ;
        RECT 14.840 32.740 16.540 34.140 ;
        RECT 16.840 32.740 18.540 34.140 ;
        RECT 18.840 32.740 20.540 34.140 ;
        RECT 20.840 32.740 22.540 34.140 ;
        RECT 22.840 32.740 24.540 34.140 ;
        RECT 24.840 32.740 26.540 34.140 ;
        RECT 26.840 32.740 28.540 34.140 ;
        RECT 28.840 32.740 30.540 34.140 ;
        RECT 30.840 32.740 32.540 34.140 ;
        RECT 32.840 32.740 34.540 34.140 ;
        RECT 34.840 32.740 36.540 34.140 ;
        RECT 36.840 32.740 38.540 34.140 ;
        RECT 38.840 32.740 40.540 34.140 ;
        RECT 40.840 32.740 42.540 34.140 ;
        RECT 42.840 32.740 44.540 34.140 ;
        RECT 44.840 32.740 46.540 34.140 ;
        RECT 46.840 32.740 48.540 34.140 ;
        RECT 48.840 32.740 50.540 34.140 ;
        RECT 50.840 32.740 52.540 34.140 ;
        RECT 52.840 32.740 54.540 34.140 ;
        RECT 54.840 32.740 56.540 34.140 ;
        RECT 56.840 32.740 58.540 34.140 ;
        RECT 58.840 32.740 60.540 34.140 ;
        RECT 60.840 32.740 62.540 34.140 ;
        RECT 62.840 32.740 64.540 34.140 ;
        RECT 64.840 32.740 66.540 34.140 ;
        RECT 66.840 32.740 68.540 34.140 ;
        RECT 68.840 32.740 70.540 34.140 ;
        RECT 70.840 32.740 72.540 34.140 ;
        RECT 72.840 32.740 74.540 34.140 ;
        RECT 86.575 32.740 88.275 34.140 ;
        RECT 88.575 32.740 90.275 34.140 ;
        RECT 90.575 32.740 92.275 34.140 ;
        RECT 92.575 32.740 94.275 34.140 ;
        RECT 94.575 32.740 96.275 34.140 ;
        RECT 96.575 32.740 98.275 34.140 ;
        RECT 98.575 32.740 100.275 34.140 ;
        RECT 100.575 32.740 102.275 34.140 ;
        RECT 102.575 32.740 104.275 34.140 ;
        RECT 104.575 32.740 106.275 34.140 ;
        RECT 106.575 32.740 108.275 34.140 ;
        RECT 108.575 32.740 110.275 34.140 ;
        RECT 110.575 32.740 112.275 34.140 ;
        RECT 112.575 32.740 114.275 34.140 ;
        RECT 114.575 32.740 116.275 34.140 ;
        RECT 116.575 32.740 118.275 34.140 ;
        RECT 118.575 32.740 120.275 34.140 ;
        RECT 120.575 32.740 122.275 34.140 ;
        RECT 122.575 32.740 124.275 34.140 ;
        RECT 124.575 32.740 126.275 34.140 ;
        RECT 126.575 32.740 128.275 34.140 ;
        RECT 128.575 32.740 130.275 34.140 ;
        RECT 130.575 32.740 132.275 34.140 ;
        RECT 132.575 32.740 134.275 34.140 ;
        RECT 134.575 32.740 136.275 34.140 ;
        RECT 136.575 32.740 138.275 34.140 ;
        RECT 138.575 32.740 140.275 34.140 ;
        RECT 140.575 32.740 142.275 34.140 ;
        RECT 142.575 32.740 144.275 34.140 ;
        RECT 144.575 32.740 146.275 34.140 ;
        RECT 146.575 32.740 148.275 34.140 ;
        RECT 148.575 32.740 150.275 34.140 ;
        RECT 150.575 32.740 152.275 34.140 ;
        RECT 152.575 32.740 154.275 34.140 ;
        RECT 6.840 30.890 8.540 32.290 ;
        RECT 8.840 30.890 10.540 32.290 ;
        RECT 10.840 30.890 12.540 32.290 ;
        RECT 12.840 30.890 14.540 32.290 ;
        RECT 14.840 30.890 16.540 32.290 ;
        RECT 16.840 30.890 18.540 32.290 ;
        RECT 18.840 30.890 20.540 32.290 ;
        RECT 20.840 30.890 22.540 32.290 ;
        RECT 22.840 30.890 24.540 32.290 ;
        RECT 24.840 30.890 26.540 32.290 ;
        RECT 26.840 30.890 28.540 32.290 ;
        RECT 28.840 30.890 30.540 32.290 ;
        RECT 30.840 30.890 32.540 32.290 ;
        RECT 32.840 30.890 34.540 32.290 ;
        RECT 34.840 30.890 36.540 32.290 ;
        RECT 36.840 30.890 38.540 32.290 ;
        RECT 38.840 30.890 40.540 32.290 ;
        RECT 40.840 30.890 42.540 32.290 ;
        RECT 42.840 30.890 44.540 32.290 ;
        RECT 44.840 30.890 46.540 32.290 ;
        RECT 46.840 30.890 48.540 32.290 ;
        RECT 48.840 30.890 50.540 32.290 ;
        RECT 50.840 30.890 52.540 32.290 ;
        RECT 52.840 30.890 54.540 32.290 ;
        RECT 54.840 30.890 56.540 32.290 ;
        RECT 56.840 30.890 58.540 32.290 ;
        RECT 58.840 30.890 60.540 32.290 ;
        RECT 60.840 30.890 62.540 32.290 ;
        RECT 62.840 30.890 64.540 32.290 ;
        RECT 64.840 30.890 66.540 32.290 ;
        RECT 66.840 30.890 68.540 32.290 ;
        RECT 68.840 30.890 70.540 32.290 ;
        RECT 70.840 30.890 72.540 32.290 ;
        RECT 72.840 30.890 74.540 32.290 ;
        RECT 86.575 30.890 88.275 32.290 ;
        RECT 88.575 30.890 90.275 32.290 ;
        RECT 90.575 30.890 92.275 32.290 ;
        RECT 92.575 30.890 94.275 32.290 ;
        RECT 94.575 30.890 96.275 32.290 ;
        RECT 96.575 30.890 98.275 32.290 ;
        RECT 98.575 30.890 100.275 32.290 ;
        RECT 100.575 30.890 102.275 32.290 ;
        RECT 102.575 30.890 104.275 32.290 ;
        RECT 104.575 30.890 106.275 32.290 ;
        RECT 106.575 30.890 108.275 32.290 ;
        RECT 108.575 30.890 110.275 32.290 ;
        RECT 110.575 30.890 112.275 32.290 ;
        RECT 112.575 30.890 114.275 32.290 ;
        RECT 114.575 30.890 116.275 32.290 ;
        RECT 116.575 30.890 118.275 32.290 ;
        RECT 118.575 30.890 120.275 32.290 ;
        RECT 120.575 30.890 122.275 32.290 ;
        RECT 122.575 30.890 124.275 32.290 ;
        RECT 124.575 30.890 126.275 32.290 ;
        RECT 126.575 30.890 128.275 32.290 ;
        RECT 128.575 30.890 130.275 32.290 ;
        RECT 130.575 30.890 132.275 32.290 ;
        RECT 132.575 30.890 134.275 32.290 ;
        RECT 134.575 30.890 136.275 32.290 ;
        RECT 136.575 30.890 138.275 32.290 ;
        RECT 138.575 30.890 140.275 32.290 ;
        RECT 140.575 30.890 142.275 32.290 ;
        RECT 142.575 30.890 144.275 32.290 ;
        RECT 144.575 30.890 146.275 32.290 ;
        RECT 146.575 30.890 148.275 32.290 ;
        RECT 148.575 30.890 150.275 32.290 ;
        RECT 150.575 30.890 152.275 32.290 ;
        RECT 152.575 30.890 154.275 32.290 ;
        RECT 6.840 29.040 8.540 30.440 ;
        RECT 8.840 29.040 10.540 30.440 ;
        RECT 10.840 29.040 12.540 30.440 ;
        RECT 12.840 29.040 14.540 30.440 ;
        RECT 14.840 29.040 16.540 30.440 ;
        RECT 16.840 29.040 18.540 30.440 ;
        RECT 18.840 29.040 20.540 30.440 ;
        RECT 20.840 29.040 22.540 30.440 ;
        RECT 22.840 29.040 24.540 30.440 ;
        RECT 24.840 29.040 26.540 30.440 ;
        RECT 26.840 29.040 28.540 30.440 ;
        RECT 28.840 29.040 30.540 30.440 ;
        RECT 30.840 29.040 32.540 30.440 ;
        RECT 32.840 29.040 34.540 30.440 ;
        RECT 34.840 29.040 36.540 30.440 ;
        RECT 36.840 29.040 38.540 30.440 ;
        RECT 38.840 29.040 40.540 30.440 ;
        RECT 40.840 29.040 42.540 30.440 ;
        RECT 42.840 29.040 44.540 30.440 ;
        RECT 44.840 29.040 46.540 30.440 ;
        RECT 46.840 29.040 48.540 30.440 ;
        RECT 48.840 29.040 50.540 30.440 ;
        RECT 50.840 29.040 52.540 30.440 ;
        RECT 52.840 29.040 54.540 30.440 ;
        RECT 54.840 29.040 56.540 30.440 ;
        RECT 56.840 29.040 58.540 30.440 ;
        RECT 58.840 29.040 60.540 30.440 ;
        RECT 60.840 29.040 62.540 30.440 ;
        RECT 62.840 29.040 64.540 30.440 ;
        RECT 64.840 29.040 66.540 30.440 ;
        RECT 66.840 29.040 68.540 30.440 ;
        RECT 68.840 29.040 70.540 30.440 ;
        RECT 70.840 29.040 72.540 30.440 ;
        RECT 72.840 29.040 74.540 30.440 ;
        RECT 86.575 29.040 88.275 30.440 ;
        RECT 88.575 29.040 90.275 30.440 ;
        RECT 90.575 29.040 92.275 30.440 ;
        RECT 92.575 29.040 94.275 30.440 ;
        RECT 94.575 29.040 96.275 30.440 ;
        RECT 96.575 29.040 98.275 30.440 ;
        RECT 98.575 29.040 100.275 30.440 ;
        RECT 100.575 29.040 102.275 30.440 ;
        RECT 102.575 29.040 104.275 30.440 ;
        RECT 104.575 29.040 106.275 30.440 ;
        RECT 106.575 29.040 108.275 30.440 ;
        RECT 108.575 29.040 110.275 30.440 ;
        RECT 110.575 29.040 112.275 30.440 ;
        RECT 112.575 29.040 114.275 30.440 ;
        RECT 114.575 29.040 116.275 30.440 ;
        RECT 116.575 29.040 118.275 30.440 ;
        RECT 118.575 29.040 120.275 30.440 ;
        RECT 120.575 29.040 122.275 30.440 ;
        RECT 122.575 29.040 124.275 30.440 ;
        RECT 124.575 29.040 126.275 30.440 ;
        RECT 126.575 29.040 128.275 30.440 ;
        RECT 128.575 29.040 130.275 30.440 ;
        RECT 130.575 29.040 132.275 30.440 ;
        RECT 132.575 29.040 134.275 30.440 ;
        RECT 134.575 29.040 136.275 30.440 ;
        RECT 136.575 29.040 138.275 30.440 ;
        RECT 138.575 29.040 140.275 30.440 ;
        RECT 140.575 29.040 142.275 30.440 ;
        RECT 142.575 29.040 144.275 30.440 ;
        RECT 144.575 29.040 146.275 30.440 ;
        RECT 146.575 29.040 148.275 30.440 ;
        RECT 148.575 29.040 150.275 30.440 ;
        RECT 150.575 29.040 152.275 30.440 ;
        RECT 152.575 29.040 154.275 30.440 ;
        RECT 6.840 27.190 8.540 28.590 ;
        RECT 8.840 27.190 10.540 28.590 ;
        RECT 10.840 27.190 12.540 28.590 ;
        RECT 12.840 27.190 14.540 28.590 ;
        RECT 14.840 27.190 16.540 28.590 ;
        RECT 16.840 27.190 18.540 28.590 ;
        RECT 18.840 27.190 20.540 28.590 ;
        RECT 20.840 27.190 22.540 28.590 ;
        RECT 22.840 27.190 24.540 28.590 ;
        RECT 24.840 27.190 26.540 28.590 ;
        RECT 26.840 27.190 28.540 28.590 ;
        RECT 28.840 27.190 30.540 28.590 ;
        RECT 30.840 27.190 32.540 28.590 ;
        RECT 32.840 27.190 34.540 28.590 ;
        RECT 34.840 27.190 36.540 28.590 ;
        RECT 36.840 27.190 38.540 28.590 ;
        RECT 38.840 27.190 40.540 28.590 ;
        RECT 40.840 27.190 42.540 28.590 ;
        RECT 42.840 27.190 44.540 28.590 ;
        RECT 44.840 27.190 46.540 28.590 ;
        RECT 46.840 27.190 48.540 28.590 ;
        RECT 48.840 27.190 50.540 28.590 ;
        RECT 50.840 27.190 52.540 28.590 ;
        RECT 52.840 27.190 54.540 28.590 ;
        RECT 54.840 27.190 56.540 28.590 ;
        RECT 56.840 27.190 58.540 28.590 ;
        RECT 58.840 27.190 60.540 28.590 ;
        RECT 60.840 27.190 62.540 28.590 ;
        RECT 62.840 27.190 64.540 28.590 ;
        RECT 64.840 27.190 66.540 28.590 ;
        RECT 66.840 27.190 68.540 28.590 ;
        RECT 68.840 27.190 70.540 28.590 ;
        RECT 70.840 27.190 72.540 28.590 ;
        RECT 72.840 27.190 74.540 28.590 ;
        RECT 86.575 27.190 88.275 28.590 ;
        RECT 88.575 27.190 90.275 28.590 ;
        RECT 90.575 27.190 92.275 28.590 ;
        RECT 92.575 27.190 94.275 28.590 ;
        RECT 94.575 27.190 96.275 28.590 ;
        RECT 96.575 27.190 98.275 28.590 ;
        RECT 98.575 27.190 100.275 28.590 ;
        RECT 100.575 27.190 102.275 28.590 ;
        RECT 102.575 27.190 104.275 28.590 ;
        RECT 104.575 27.190 106.275 28.590 ;
        RECT 106.575 27.190 108.275 28.590 ;
        RECT 108.575 27.190 110.275 28.590 ;
        RECT 110.575 27.190 112.275 28.590 ;
        RECT 112.575 27.190 114.275 28.590 ;
        RECT 114.575 27.190 116.275 28.590 ;
        RECT 116.575 27.190 118.275 28.590 ;
        RECT 118.575 27.190 120.275 28.590 ;
        RECT 120.575 27.190 122.275 28.590 ;
        RECT 122.575 27.190 124.275 28.590 ;
        RECT 124.575 27.190 126.275 28.590 ;
        RECT 126.575 27.190 128.275 28.590 ;
        RECT 128.575 27.190 130.275 28.590 ;
        RECT 130.575 27.190 132.275 28.590 ;
        RECT 132.575 27.190 134.275 28.590 ;
        RECT 134.575 27.190 136.275 28.590 ;
        RECT 136.575 27.190 138.275 28.590 ;
        RECT 138.575 27.190 140.275 28.590 ;
        RECT 140.575 27.190 142.275 28.590 ;
        RECT 142.575 27.190 144.275 28.590 ;
        RECT 144.575 27.190 146.275 28.590 ;
        RECT 146.575 27.190 148.275 28.590 ;
        RECT 148.575 27.190 150.275 28.590 ;
        RECT 150.575 27.190 152.275 28.590 ;
        RECT 152.575 27.190 154.275 28.590 ;
        RECT 6.840 25.340 8.540 26.740 ;
        RECT 8.840 25.340 10.540 26.740 ;
        RECT 10.840 25.340 12.540 26.740 ;
        RECT 12.840 25.340 14.540 26.740 ;
        RECT 14.840 25.340 16.540 26.740 ;
        RECT 16.840 25.340 18.540 26.740 ;
        RECT 18.840 25.340 20.540 26.740 ;
        RECT 20.840 25.340 22.540 26.740 ;
        RECT 22.840 25.340 24.540 26.740 ;
        RECT 24.840 25.340 26.540 26.740 ;
        RECT 26.840 25.340 28.540 26.740 ;
        RECT 28.840 25.340 30.540 26.740 ;
        RECT 30.840 25.340 32.540 26.740 ;
        RECT 32.840 25.340 34.540 26.740 ;
        RECT 34.840 25.340 36.540 26.740 ;
        RECT 36.840 25.340 38.540 26.740 ;
        RECT 38.840 25.340 40.540 26.740 ;
        RECT 40.840 25.340 42.540 26.740 ;
        RECT 42.840 25.340 44.540 26.740 ;
        RECT 44.840 25.340 46.540 26.740 ;
        RECT 46.840 25.340 48.540 26.740 ;
        RECT 48.840 25.340 50.540 26.740 ;
        RECT 50.840 25.340 52.540 26.740 ;
        RECT 52.840 25.340 54.540 26.740 ;
        RECT 54.840 25.340 56.540 26.740 ;
        RECT 56.840 25.340 58.540 26.740 ;
        RECT 58.840 25.340 60.540 26.740 ;
        RECT 60.840 25.340 62.540 26.740 ;
        RECT 62.840 25.340 64.540 26.740 ;
        RECT 64.840 25.340 66.540 26.740 ;
        RECT 66.840 25.340 68.540 26.740 ;
        RECT 68.840 25.340 70.540 26.740 ;
        RECT 70.840 25.340 72.540 26.740 ;
        RECT 72.840 25.340 74.540 26.740 ;
        RECT 86.575 25.340 88.275 26.740 ;
        RECT 88.575 25.340 90.275 26.740 ;
        RECT 90.575 25.340 92.275 26.740 ;
        RECT 92.575 25.340 94.275 26.740 ;
        RECT 94.575 25.340 96.275 26.740 ;
        RECT 96.575 25.340 98.275 26.740 ;
        RECT 98.575 25.340 100.275 26.740 ;
        RECT 100.575 25.340 102.275 26.740 ;
        RECT 102.575 25.340 104.275 26.740 ;
        RECT 104.575 25.340 106.275 26.740 ;
        RECT 106.575 25.340 108.275 26.740 ;
        RECT 108.575 25.340 110.275 26.740 ;
        RECT 110.575 25.340 112.275 26.740 ;
        RECT 112.575 25.340 114.275 26.740 ;
        RECT 114.575 25.340 116.275 26.740 ;
        RECT 116.575 25.340 118.275 26.740 ;
        RECT 118.575 25.340 120.275 26.740 ;
        RECT 120.575 25.340 122.275 26.740 ;
        RECT 122.575 25.340 124.275 26.740 ;
        RECT 124.575 25.340 126.275 26.740 ;
        RECT 126.575 25.340 128.275 26.740 ;
        RECT 128.575 25.340 130.275 26.740 ;
        RECT 130.575 25.340 132.275 26.740 ;
        RECT 132.575 25.340 134.275 26.740 ;
        RECT 134.575 25.340 136.275 26.740 ;
        RECT 136.575 25.340 138.275 26.740 ;
        RECT 138.575 25.340 140.275 26.740 ;
        RECT 140.575 25.340 142.275 26.740 ;
        RECT 142.575 25.340 144.275 26.740 ;
        RECT 144.575 25.340 146.275 26.740 ;
        RECT 146.575 25.340 148.275 26.740 ;
        RECT 148.575 25.340 150.275 26.740 ;
        RECT 150.575 25.340 152.275 26.740 ;
        RECT 152.575 25.340 154.275 26.740 ;
        RECT 6.840 23.490 8.540 24.890 ;
        RECT 8.840 23.490 10.540 24.890 ;
        RECT 10.840 23.490 12.540 24.890 ;
        RECT 12.840 23.490 14.540 24.890 ;
        RECT 14.840 23.490 16.540 24.890 ;
        RECT 16.840 23.490 18.540 24.890 ;
        RECT 18.840 23.490 20.540 24.890 ;
        RECT 20.840 23.490 22.540 24.890 ;
        RECT 22.840 23.490 24.540 24.890 ;
        RECT 24.840 23.490 26.540 24.890 ;
        RECT 26.840 23.490 28.540 24.890 ;
        RECT 28.840 23.490 30.540 24.890 ;
        RECT 30.840 23.490 32.540 24.890 ;
        RECT 32.840 23.490 34.540 24.890 ;
        RECT 34.840 23.490 36.540 24.890 ;
        RECT 36.840 23.490 38.540 24.890 ;
        RECT 38.840 23.490 40.540 24.890 ;
        RECT 40.840 23.490 42.540 24.890 ;
        RECT 42.840 23.490 44.540 24.890 ;
        RECT 44.840 23.490 46.540 24.890 ;
        RECT 46.840 23.490 48.540 24.890 ;
        RECT 48.840 23.490 50.540 24.890 ;
        RECT 50.840 23.490 52.540 24.890 ;
        RECT 52.840 23.490 54.540 24.890 ;
        RECT 54.840 23.490 56.540 24.890 ;
        RECT 56.840 23.490 58.540 24.890 ;
        RECT 58.840 23.490 60.540 24.890 ;
        RECT 60.840 23.490 62.540 24.890 ;
        RECT 62.840 23.490 64.540 24.890 ;
        RECT 64.840 23.490 66.540 24.890 ;
        RECT 66.840 23.490 68.540 24.890 ;
        RECT 68.840 23.490 70.540 24.890 ;
        RECT 70.840 23.490 72.540 24.890 ;
        RECT 72.840 23.490 74.540 24.890 ;
        RECT 86.575 23.490 88.275 24.890 ;
        RECT 88.575 23.490 90.275 24.890 ;
        RECT 90.575 23.490 92.275 24.890 ;
        RECT 92.575 23.490 94.275 24.890 ;
        RECT 94.575 23.490 96.275 24.890 ;
        RECT 96.575 23.490 98.275 24.890 ;
        RECT 98.575 23.490 100.275 24.890 ;
        RECT 100.575 23.490 102.275 24.890 ;
        RECT 102.575 23.490 104.275 24.890 ;
        RECT 104.575 23.490 106.275 24.890 ;
        RECT 106.575 23.490 108.275 24.890 ;
        RECT 108.575 23.490 110.275 24.890 ;
        RECT 110.575 23.490 112.275 24.890 ;
        RECT 112.575 23.490 114.275 24.890 ;
        RECT 114.575 23.490 116.275 24.890 ;
        RECT 116.575 23.490 118.275 24.890 ;
        RECT 118.575 23.490 120.275 24.890 ;
        RECT 120.575 23.490 122.275 24.890 ;
        RECT 122.575 23.490 124.275 24.890 ;
        RECT 124.575 23.490 126.275 24.890 ;
        RECT 126.575 23.490 128.275 24.890 ;
        RECT 128.575 23.490 130.275 24.890 ;
        RECT 130.575 23.490 132.275 24.890 ;
        RECT 132.575 23.490 134.275 24.890 ;
        RECT 134.575 23.490 136.275 24.890 ;
        RECT 136.575 23.490 138.275 24.890 ;
        RECT 138.575 23.490 140.275 24.890 ;
        RECT 140.575 23.490 142.275 24.890 ;
        RECT 142.575 23.490 144.275 24.890 ;
        RECT 144.575 23.490 146.275 24.890 ;
        RECT 146.575 23.490 148.275 24.890 ;
        RECT 148.575 23.490 150.275 24.890 ;
        RECT 150.575 23.490 152.275 24.890 ;
        RECT 152.575 23.490 154.275 24.890 ;
        RECT 6.840 21.640 8.540 23.040 ;
        RECT 8.840 21.640 10.540 23.040 ;
        RECT 10.840 21.640 12.540 23.040 ;
        RECT 12.840 21.640 14.540 23.040 ;
        RECT 14.840 21.640 16.540 23.040 ;
        RECT 16.840 21.640 18.540 23.040 ;
        RECT 18.840 21.640 20.540 23.040 ;
        RECT 20.840 21.640 22.540 23.040 ;
        RECT 22.840 21.640 24.540 23.040 ;
        RECT 24.840 21.640 26.540 23.040 ;
        RECT 26.840 21.640 28.540 23.040 ;
        RECT 28.840 21.640 30.540 23.040 ;
        RECT 30.840 21.640 32.540 23.040 ;
        RECT 32.840 21.640 34.540 23.040 ;
        RECT 34.840 21.640 36.540 23.040 ;
        RECT 36.840 21.640 38.540 23.040 ;
        RECT 38.840 21.640 40.540 23.040 ;
        RECT 40.840 21.640 42.540 23.040 ;
        RECT 42.840 21.640 44.540 23.040 ;
        RECT 44.840 21.640 46.540 23.040 ;
        RECT 46.840 21.640 48.540 23.040 ;
        RECT 48.840 21.640 50.540 23.040 ;
        RECT 50.840 21.640 52.540 23.040 ;
        RECT 52.840 21.640 54.540 23.040 ;
        RECT 54.840 21.640 56.540 23.040 ;
        RECT 56.840 21.640 58.540 23.040 ;
        RECT 58.840 21.640 60.540 23.040 ;
        RECT 60.840 21.640 62.540 23.040 ;
        RECT 62.840 21.640 64.540 23.040 ;
        RECT 64.840 21.640 66.540 23.040 ;
        RECT 66.840 21.640 68.540 23.040 ;
        RECT 68.840 21.640 70.540 23.040 ;
        RECT 70.840 21.640 72.540 23.040 ;
        RECT 72.840 21.640 74.540 23.040 ;
        RECT 86.575 21.640 88.275 23.040 ;
        RECT 88.575 21.640 90.275 23.040 ;
        RECT 90.575 21.640 92.275 23.040 ;
        RECT 92.575 21.640 94.275 23.040 ;
        RECT 94.575 21.640 96.275 23.040 ;
        RECT 96.575 21.640 98.275 23.040 ;
        RECT 98.575 21.640 100.275 23.040 ;
        RECT 100.575 21.640 102.275 23.040 ;
        RECT 102.575 21.640 104.275 23.040 ;
        RECT 104.575 21.640 106.275 23.040 ;
        RECT 106.575 21.640 108.275 23.040 ;
        RECT 108.575 21.640 110.275 23.040 ;
        RECT 110.575 21.640 112.275 23.040 ;
        RECT 112.575 21.640 114.275 23.040 ;
        RECT 114.575 21.640 116.275 23.040 ;
        RECT 116.575 21.640 118.275 23.040 ;
        RECT 118.575 21.640 120.275 23.040 ;
        RECT 120.575 21.640 122.275 23.040 ;
        RECT 122.575 21.640 124.275 23.040 ;
        RECT 124.575 21.640 126.275 23.040 ;
        RECT 126.575 21.640 128.275 23.040 ;
        RECT 128.575 21.640 130.275 23.040 ;
        RECT 130.575 21.640 132.275 23.040 ;
        RECT 132.575 21.640 134.275 23.040 ;
        RECT 134.575 21.640 136.275 23.040 ;
        RECT 136.575 21.640 138.275 23.040 ;
        RECT 138.575 21.640 140.275 23.040 ;
        RECT 140.575 21.640 142.275 23.040 ;
        RECT 142.575 21.640 144.275 23.040 ;
        RECT 144.575 21.640 146.275 23.040 ;
        RECT 146.575 21.640 148.275 23.040 ;
        RECT 148.575 21.640 150.275 23.040 ;
        RECT 150.575 21.640 152.275 23.040 ;
        RECT 152.575 21.640 154.275 23.040 ;
        RECT 6.840 19.790 8.540 21.190 ;
        RECT 8.840 19.790 10.540 21.190 ;
        RECT 10.840 19.790 12.540 21.190 ;
        RECT 12.840 19.790 14.540 21.190 ;
        RECT 14.840 19.790 16.540 21.190 ;
        RECT 16.840 19.790 18.540 21.190 ;
        RECT 18.840 19.790 20.540 21.190 ;
        RECT 20.840 19.790 22.540 21.190 ;
        RECT 22.840 19.790 24.540 21.190 ;
        RECT 24.840 19.790 26.540 21.190 ;
        RECT 26.840 19.790 28.540 21.190 ;
        RECT 28.840 19.790 30.540 21.190 ;
        RECT 30.840 19.790 32.540 21.190 ;
        RECT 32.840 19.790 34.540 21.190 ;
        RECT 34.840 19.790 36.540 21.190 ;
        RECT 36.840 19.790 38.540 21.190 ;
        RECT 38.840 19.790 40.540 21.190 ;
        RECT 40.840 19.790 42.540 21.190 ;
        RECT 42.840 19.790 44.540 21.190 ;
        RECT 44.840 19.790 46.540 21.190 ;
        RECT 46.840 19.790 48.540 21.190 ;
        RECT 48.840 19.790 50.540 21.190 ;
        RECT 50.840 19.790 52.540 21.190 ;
        RECT 52.840 19.790 54.540 21.190 ;
        RECT 54.840 19.790 56.540 21.190 ;
        RECT 56.840 19.790 58.540 21.190 ;
        RECT 58.840 19.790 60.540 21.190 ;
        RECT 60.840 19.790 62.540 21.190 ;
        RECT 62.840 19.790 64.540 21.190 ;
        RECT 64.840 19.790 66.540 21.190 ;
        RECT 66.840 19.790 68.540 21.190 ;
        RECT 68.840 19.790 70.540 21.190 ;
        RECT 70.840 19.790 72.540 21.190 ;
        RECT 72.840 19.790 74.540 21.190 ;
        RECT 86.575 19.790 88.275 21.190 ;
        RECT 88.575 19.790 90.275 21.190 ;
        RECT 90.575 19.790 92.275 21.190 ;
        RECT 92.575 19.790 94.275 21.190 ;
        RECT 94.575 19.790 96.275 21.190 ;
        RECT 96.575 19.790 98.275 21.190 ;
        RECT 98.575 19.790 100.275 21.190 ;
        RECT 100.575 19.790 102.275 21.190 ;
        RECT 102.575 19.790 104.275 21.190 ;
        RECT 104.575 19.790 106.275 21.190 ;
        RECT 106.575 19.790 108.275 21.190 ;
        RECT 108.575 19.790 110.275 21.190 ;
        RECT 110.575 19.790 112.275 21.190 ;
        RECT 112.575 19.790 114.275 21.190 ;
        RECT 114.575 19.790 116.275 21.190 ;
        RECT 116.575 19.790 118.275 21.190 ;
        RECT 118.575 19.790 120.275 21.190 ;
        RECT 120.575 19.790 122.275 21.190 ;
        RECT 122.575 19.790 124.275 21.190 ;
        RECT 124.575 19.790 126.275 21.190 ;
        RECT 126.575 19.790 128.275 21.190 ;
        RECT 128.575 19.790 130.275 21.190 ;
        RECT 130.575 19.790 132.275 21.190 ;
        RECT 132.575 19.790 134.275 21.190 ;
        RECT 134.575 19.790 136.275 21.190 ;
        RECT 136.575 19.790 138.275 21.190 ;
        RECT 138.575 19.790 140.275 21.190 ;
        RECT 140.575 19.790 142.275 21.190 ;
        RECT 142.575 19.790 144.275 21.190 ;
        RECT 144.575 19.790 146.275 21.190 ;
        RECT 146.575 19.790 148.275 21.190 ;
        RECT 148.575 19.790 150.275 21.190 ;
        RECT 150.575 19.790 152.275 21.190 ;
        RECT 152.575 19.790 154.275 21.190 ;
        RECT 6.840 17.940 8.540 19.340 ;
        RECT 8.840 17.940 10.540 19.340 ;
        RECT 10.840 17.940 12.540 19.340 ;
        RECT 12.840 17.940 14.540 19.340 ;
        RECT 14.840 17.940 16.540 19.340 ;
        RECT 16.840 17.940 18.540 19.340 ;
        RECT 18.840 17.940 20.540 19.340 ;
        RECT 20.840 17.940 22.540 19.340 ;
        RECT 22.840 17.940 24.540 19.340 ;
        RECT 24.840 17.940 26.540 19.340 ;
        RECT 26.840 17.940 28.540 19.340 ;
        RECT 28.840 17.940 30.540 19.340 ;
        RECT 30.840 17.940 32.540 19.340 ;
        RECT 32.840 17.940 34.540 19.340 ;
        RECT 34.840 17.940 36.540 19.340 ;
        RECT 36.840 17.940 38.540 19.340 ;
        RECT 38.840 17.940 40.540 19.340 ;
        RECT 40.840 17.940 42.540 19.340 ;
        RECT 42.840 17.940 44.540 19.340 ;
        RECT 44.840 17.940 46.540 19.340 ;
        RECT 46.840 17.940 48.540 19.340 ;
        RECT 48.840 17.940 50.540 19.340 ;
        RECT 50.840 17.940 52.540 19.340 ;
        RECT 52.840 17.940 54.540 19.340 ;
        RECT 54.840 17.940 56.540 19.340 ;
        RECT 56.840 17.940 58.540 19.340 ;
        RECT 58.840 17.940 60.540 19.340 ;
        RECT 60.840 17.940 62.540 19.340 ;
        RECT 62.840 17.940 64.540 19.340 ;
        RECT 64.840 17.940 66.540 19.340 ;
        RECT 66.840 17.940 68.540 19.340 ;
        RECT 68.840 17.940 70.540 19.340 ;
        RECT 70.840 17.940 72.540 19.340 ;
        RECT 72.840 17.940 74.540 19.340 ;
        RECT 86.575 17.940 88.275 19.340 ;
        RECT 88.575 17.940 90.275 19.340 ;
        RECT 90.575 17.940 92.275 19.340 ;
        RECT 92.575 17.940 94.275 19.340 ;
        RECT 94.575 17.940 96.275 19.340 ;
        RECT 96.575 17.940 98.275 19.340 ;
        RECT 98.575 17.940 100.275 19.340 ;
        RECT 100.575 17.940 102.275 19.340 ;
        RECT 102.575 17.940 104.275 19.340 ;
        RECT 104.575 17.940 106.275 19.340 ;
        RECT 106.575 17.940 108.275 19.340 ;
        RECT 108.575 17.940 110.275 19.340 ;
        RECT 110.575 17.940 112.275 19.340 ;
        RECT 112.575 17.940 114.275 19.340 ;
        RECT 114.575 17.940 116.275 19.340 ;
        RECT 116.575 17.940 118.275 19.340 ;
        RECT 118.575 17.940 120.275 19.340 ;
        RECT 120.575 17.940 122.275 19.340 ;
        RECT 122.575 17.940 124.275 19.340 ;
        RECT 124.575 17.940 126.275 19.340 ;
        RECT 126.575 17.940 128.275 19.340 ;
        RECT 128.575 17.940 130.275 19.340 ;
        RECT 130.575 17.940 132.275 19.340 ;
        RECT 132.575 17.940 134.275 19.340 ;
        RECT 134.575 17.940 136.275 19.340 ;
        RECT 136.575 17.940 138.275 19.340 ;
        RECT 138.575 17.940 140.275 19.340 ;
        RECT 140.575 17.940 142.275 19.340 ;
        RECT 142.575 17.940 144.275 19.340 ;
        RECT 144.575 17.940 146.275 19.340 ;
        RECT 146.575 17.940 148.275 19.340 ;
        RECT 148.575 17.940 150.275 19.340 ;
        RECT 150.575 17.940 152.275 19.340 ;
        RECT 152.575 17.940 154.275 19.340 ;
        RECT 6.840 16.090 8.540 17.490 ;
        RECT 8.840 16.090 10.540 17.490 ;
        RECT 10.840 16.090 12.540 17.490 ;
        RECT 12.840 16.090 14.540 17.490 ;
        RECT 14.840 16.090 16.540 17.490 ;
        RECT 16.840 16.090 18.540 17.490 ;
        RECT 18.840 16.090 20.540 17.490 ;
        RECT 20.840 16.090 22.540 17.490 ;
        RECT 22.840 16.090 24.540 17.490 ;
        RECT 24.840 16.090 26.540 17.490 ;
        RECT 26.840 16.090 28.540 17.490 ;
        RECT 28.840 16.090 30.540 17.490 ;
        RECT 30.840 16.090 32.540 17.490 ;
        RECT 32.840 16.090 34.540 17.490 ;
        RECT 34.840 16.090 36.540 17.490 ;
        RECT 36.840 16.090 38.540 17.490 ;
        RECT 38.840 16.090 40.540 17.490 ;
        RECT 40.840 16.090 42.540 17.490 ;
        RECT 42.840 16.090 44.540 17.490 ;
        RECT 44.840 16.090 46.540 17.490 ;
        RECT 46.840 16.090 48.540 17.490 ;
        RECT 48.840 16.090 50.540 17.490 ;
        RECT 50.840 16.090 52.540 17.490 ;
        RECT 52.840 16.090 54.540 17.490 ;
        RECT 54.840 16.090 56.540 17.490 ;
        RECT 56.840 16.090 58.540 17.490 ;
        RECT 58.840 16.090 60.540 17.490 ;
        RECT 60.840 16.090 62.540 17.490 ;
        RECT 62.840 16.090 64.540 17.490 ;
        RECT 64.840 16.090 66.540 17.490 ;
        RECT 66.840 16.090 68.540 17.490 ;
        RECT 68.840 16.090 70.540 17.490 ;
        RECT 70.840 16.090 72.540 17.490 ;
        RECT 72.840 16.090 74.540 17.490 ;
        RECT 86.575 16.090 88.275 17.490 ;
        RECT 88.575 16.090 90.275 17.490 ;
        RECT 90.575 16.090 92.275 17.490 ;
        RECT 92.575 16.090 94.275 17.490 ;
        RECT 94.575 16.090 96.275 17.490 ;
        RECT 96.575 16.090 98.275 17.490 ;
        RECT 98.575 16.090 100.275 17.490 ;
        RECT 100.575 16.090 102.275 17.490 ;
        RECT 102.575 16.090 104.275 17.490 ;
        RECT 104.575 16.090 106.275 17.490 ;
        RECT 106.575 16.090 108.275 17.490 ;
        RECT 108.575 16.090 110.275 17.490 ;
        RECT 110.575 16.090 112.275 17.490 ;
        RECT 112.575 16.090 114.275 17.490 ;
        RECT 114.575 16.090 116.275 17.490 ;
        RECT 116.575 16.090 118.275 17.490 ;
        RECT 118.575 16.090 120.275 17.490 ;
        RECT 120.575 16.090 122.275 17.490 ;
        RECT 122.575 16.090 124.275 17.490 ;
        RECT 124.575 16.090 126.275 17.490 ;
        RECT 126.575 16.090 128.275 17.490 ;
        RECT 128.575 16.090 130.275 17.490 ;
        RECT 130.575 16.090 132.275 17.490 ;
        RECT 132.575 16.090 134.275 17.490 ;
        RECT 134.575 16.090 136.275 17.490 ;
        RECT 136.575 16.090 138.275 17.490 ;
        RECT 138.575 16.090 140.275 17.490 ;
        RECT 140.575 16.090 142.275 17.490 ;
        RECT 142.575 16.090 144.275 17.490 ;
        RECT 144.575 16.090 146.275 17.490 ;
        RECT 146.575 16.090 148.275 17.490 ;
        RECT 148.575 16.090 150.275 17.490 ;
        RECT 150.575 16.090 152.275 17.490 ;
        RECT 152.575 16.090 154.275 17.490 ;
        RECT 6.840 14.240 8.540 15.640 ;
        RECT 8.840 14.240 10.540 15.640 ;
        RECT 10.840 14.240 12.540 15.640 ;
        RECT 12.840 14.240 14.540 15.640 ;
        RECT 14.840 14.240 16.540 15.640 ;
        RECT 16.840 14.240 18.540 15.640 ;
        RECT 18.840 14.240 20.540 15.640 ;
        RECT 20.840 14.240 22.540 15.640 ;
        RECT 22.840 14.240 24.540 15.640 ;
        RECT 24.840 14.240 26.540 15.640 ;
        RECT 26.840 14.240 28.540 15.640 ;
        RECT 28.840 14.240 30.540 15.640 ;
        RECT 30.840 14.240 32.540 15.640 ;
        RECT 32.840 14.240 34.540 15.640 ;
        RECT 34.840 14.240 36.540 15.640 ;
        RECT 36.840 14.240 38.540 15.640 ;
        RECT 38.840 14.240 40.540 15.640 ;
        RECT 40.840 14.240 42.540 15.640 ;
        RECT 42.840 14.240 44.540 15.640 ;
        RECT 44.840 14.240 46.540 15.640 ;
        RECT 46.840 14.240 48.540 15.640 ;
        RECT 48.840 14.240 50.540 15.640 ;
        RECT 50.840 14.240 52.540 15.640 ;
        RECT 52.840 14.240 54.540 15.640 ;
        RECT 54.840 14.240 56.540 15.640 ;
        RECT 56.840 14.240 58.540 15.640 ;
        RECT 58.840 14.240 60.540 15.640 ;
        RECT 60.840 14.240 62.540 15.640 ;
        RECT 62.840 14.240 64.540 15.640 ;
        RECT 64.840 14.240 66.540 15.640 ;
        RECT 66.840 14.240 68.540 15.640 ;
        RECT 68.840 14.240 70.540 15.640 ;
        RECT 70.840 14.240 72.540 15.640 ;
        RECT 72.840 14.240 74.540 15.640 ;
        RECT 86.575 14.240 88.275 15.640 ;
        RECT 88.575 14.240 90.275 15.640 ;
        RECT 90.575 14.240 92.275 15.640 ;
        RECT 92.575 14.240 94.275 15.640 ;
        RECT 94.575 14.240 96.275 15.640 ;
        RECT 96.575 14.240 98.275 15.640 ;
        RECT 98.575 14.240 100.275 15.640 ;
        RECT 100.575 14.240 102.275 15.640 ;
        RECT 102.575 14.240 104.275 15.640 ;
        RECT 104.575 14.240 106.275 15.640 ;
        RECT 106.575 14.240 108.275 15.640 ;
        RECT 108.575 14.240 110.275 15.640 ;
        RECT 110.575 14.240 112.275 15.640 ;
        RECT 112.575 14.240 114.275 15.640 ;
        RECT 114.575 14.240 116.275 15.640 ;
        RECT 116.575 14.240 118.275 15.640 ;
        RECT 118.575 14.240 120.275 15.640 ;
        RECT 120.575 14.240 122.275 15.640 ;
        RECT 122.575 14.240 124.275 15.640 ;
        RECT 124.575 14.240 126.275 15.640 ;
        RECT 126.575 14.240 128.275 15.640 ;
        RECT 128.575 14.240 130.275 15.640 ;
        RECT 130.575 14.240 132.275 15.640 ;
        RECT 132.575 14.240 134.275 15.640 ;
        RECT 134.575 14.240 136.275 15.640 ;
        RECT 136.575 14.240 138.275 15.640 ;
        RECT 138.575 14.240 140.275 15.640 ;
        RECT 140.575 14.240 142.275 15.640 ;
        RECT 142.575 14.240 144.275 15.640 ;
        RECT 144.575 14.240 146.275 15.640 ;
        RECT 146.575 14.240 148.275 15.640 ;
        RECT 148.575 14.240 150.275 15.640 ;
        RECT 150.575 14.240 152.275 15.640 ;
        RECT 152.575 14.240 154.275 15.640 ;
        RECT 6.840 12.390 8.540 13.790 ;
        RECT 8.840 12.390 10.540 13.790 ;
        RECT 10.840 12.390 12.540 13.790 ;
        RECT 12.840 12.390 14.540 13.790 ;
        RECT 14.840 12.390 16.540 13.790 ;
        RECT 16.840 12.390 18.540 13.790 ;
        RECT 18.840 12.390 20.540 13.790 ;
        RECT 20.840 12.390 22.540 13.790 ;
        RECT 22.840 12.390 24.540 13.790 ;
        RECT 24.840 12.390 26.540 13.790 ;
        RECT 26.840 12.390 28.540 13.790 ;
        RECT 28.840 12.390 30.540 13.790 ;
        RECT 30.840 12.390 32.540 13.790 ;
        RECT 32.840 12.390 34.540 13.790 ;
        RECT 34.840 12.390 36.540 13.790 ;
        RECT 36.840 12.390 38.540 13.790 ;
        RECT 38.840 12.390 40.540 13.790 ;
        RECT 40.840 12.390 42.540 13.790 ;
        RECT 42.840 12.390 44.540 13.790 ;
        RECT 44.840 12.390 46.540 13.790 ;
        RECT 46.840 12.390 48.540 13.790 ;
        RECT 48.840 12.390 50.540 13.790 ;
        RECT 50.840 12.390 52.540 13.790 ;
        RECT 52.840 12.390 54.540 13.790 ;
        RECT 54.840 12.390 56.540 13.790 ;
        RECT 56.840 12.390 58.540 13.790 ;
        RECT 58.840 12.390 60.540 13.790 ;
        RECT 60.840 12.390 62.540 13.790 ;
        RECT 62.840 12.390 64.540 13.790 ;
        RECT 64.840 12.390 66.540 13.790 ;
        RECT 66.840 12.390 68.540 13.790 ;
        RECT 68.840 12.390 70.540 13.790 ;
        RECT 70.840 12.390 72.540 13.790 ;
        RECT 72.840 12.390 74.540 13.790 ;
        RECT 86.575 12.390 88.275 13.790 ;
        RECT 88.575 12.390 90.275 13.790 ;
        RECT 90.575 12.390 92.275 13.790 ;
        RECT 92.575 12.390 94.275 13.790 ;
        RECT 94.575 12.390 96.275 13.790 ;
        RECT 96.575 12.390 98.275 13.790 ;
        RECT 98.575 12.390 100.275 13.790 ;
        RECT 100.575 12.390 102.275 13.790 ;
        RECT 102.575 12.390 104.275 13.790 ;
        RECT 104.575 12.390 106.275 13.790 ;
        RECT 106.575 12.390 108.275 13.790 ;
        RECT 108.575 12.390 110.275 13.790 ;
        RECT 110.575 12.390 112.275 13.790 ;
        RECT 112.575 12.390 114.275 13.790 ;
        RECT 114.575 12.390 116.275 13.790 ;
        RECT 116.575 12.390 118.275 13.790 ;
        RECT 118.575 12.390 120.275 13.790 ;
        RECT 120.575 12.390 122.275 13.790 ;
        RECT 122.575 12.390 124.275 13.790 ;
        RECT 124.575 12.390 126.275 13.790 ;
        RECT 126.575 12.390 128.275 13.790 ;
        RECT 128.575 12.390 130.275 13.790 ;
        RECT 130.575 12.390 132.275 13.790 ;
        RECT 132.575 12.390 134.275 13.790 ;
        RECT 134.575 12.390 136.275 13.790 ;
        RECT 136.575 12.390 138.275 13.790 ;
        RECT 138.575 12.390 140.275 13.790 ;
        RECT 140.575 12.390 142.275 13.790 ;
        RECT 142.575 12.390 144.275 13.790 ;
        RECT 144.575 12.390 146.275 13.790 ;
        RECT 146.575 12.390 148.275 13.790 ;
        RECT 148.575 12.390 150.275 13.790 ;
        RECT 150.575 12.390 152.275 13.790 ;
        RECT 152.575 12.390 154.275 13.790 ;
        RECT 6.840 10.540 8.540 11.940 ;
        RECT 8.840 10.540 10.540 11.940 ;
        RECT 10.840 10.540 12.540 11.940 ;
        RECT 12.840 10.540 14.540 11.940 ;
        RECT 14.840 10.540 16.540 11.940 ;
        RECT 16.840 10.540 18.540 11.940 ;
        RECT 18.840 10.540 20.540 11.940 ;
        RECT 20.840 10.540 22.540 11.940 ;
        RECT 22.840 10.540 24.540 11.940 ;
        RECT 24.840 10.540 26.540 11.940 ;
        RECT 26.840 10.540 28.540 11.940 ;
        RECT 28.840 10.540 30.540 11.940 ;
        RECT 30.840 10.540 32.540 11.940 ;
        RECT 32.840 10.540 34.540 11.940 ;
        RECT 34.840 10.540 36.540 11.940 ;
        RECT 36.840 10.540 38.540 11.940 ;
        RECT 38.840 10.540 40.540 11.940 ;
        RECT 40.840 10.540 42.540 11.940 ;
        RECT 42.840 10.540 44.540 11.940 ;
        RECT 44.840 10.540 46.540 11.940 ;
        RECT 46.840 10.540 48.540 11.940 ;
        RECT 48.840 10.540 50.540 11.940 ;
        RECT 50.840 10.540 52.540 11.940 ;
        RECT 52.840 10.540 54.540 11.940 ;
        RECT 54.840 10.540 56.540 11.940 ;
        RECT 56.840 10.540 58.540 11.940 ;
        RECT 58.840 10.540 60.540 11.940 ;
        RECT 60.840 10.540 62.540 11.940 ;
        RECT 62.840 10.540 64.540 11.940 ;
        RECT 64.840 10.540 66.540 11.940 ;
        RECT 66.840 10.540 68.540 11.940 ;
        RECT 68.840 10.540 70.540 11.940 ;
        RECT 70.840 10.540 72.540 11.940 ;
        RECT 72.840 10.540 74.540 11.940 ;
        RECT 86.575 10.540 88.275 11.940 ;
        RECT 88.575 10.540 90.275 11.940 ;
        RECT 90.575 10.540 92.275 11.940 ;
        RECT 92.575 10.540 94.275 11.940 ;
        RECT 94.575 10.540 96.275 11.940 ;
        RECT 96.575 10.540 98.275 11.940 ;
        RECT 98.575 10.540 100.275 11.940 ;
        RECT 100.575 10.540 102.275 11.940 ;
        RECT 102.575 10.540 104.275 11.940 ;
        RECT 104.575 10.540 106.275 11.940 ;
        RECT 106.575 10.540 108.275 11.940 ;
        RECT 108.575 10.540 110.275 11.940 ;
        RECT 110.575 10.540 112.275 11.940 ;
        RECT 112.575 10.540 114.275 11.940 ;
        RECT 114.575 10.540 116.275 11.940 ;
        RECT 116.575 10.540 118.275 11.940 ;
        RECT 118.575 10.540 120.275 11.940 ;
        RECT 120.575 10.540 122.275 11.940 ;
        RECT 122.575 10.540 124.275 11.940 ;
        RECT 124.575 10.540 126.275 11.940 ;
        RECT 126.575 10.540 128.275 11.940 ;
        RECT 128.575 10.540 130.275 11.940 ;
        RECT 130.575 10.540 132.275 11.940 ;
        RECT 132.575 10.540 134.275 11.940 ;
        RECT 134.575 10.540 136.275 11.940 ;
        RECT 136.575 10.540 138.275 11.940 ;
        RECT 138.575 10.540 140.275 11.940 ;
        RECT 140.575 10.540 142.275 11.940 ;
        RECT 142.575 10.540 144.275 11.940 ;
        RECT 144.575 10.540 146.275 11.940 ;
        RECT 146.575 10.540 148.275 11.940 ;
        RECT 148.575 10.540 150.275 11.940 ;
        RECT 150.575 10.540 152.275 11.940 ;
        RECT 152.575 10.540 154.275 11.940 ;
        RECT 6.840 8.690 8.540 10.090 ;
        RECT 8.840 8.690 10.540 10.090 ;
        RECT 10.840 8.690 12.540 10.090 ;
        RECT 12.840 8.690 14.540 10.090 ;
        RECT 14.840 8.690 16.540 10.090 ;
        RECT 16.840 8.690 18.540 10.090 ;
        RECT 18.840 8.690 20.540 10.090 ;
        RECT 20.840 8.690 22.540 10.090 ;
        RECT 22.840 8.690 24.540 10.090 ;
        RECT 24.840 8.690 26.540 10.090 ;
        RECT 26.840 8.690 28.540 10.090 ;
        RECT 28.840 8.690 30.540 10.090 ;
        RECT 30.840 8.690 32.540 10.090 ;
        RECT 32.840 8.690 34.540 10.090 ;
        RECT 34.840 8.690 36.540 10.090 ;
        RECT 36.840 8.690 38.540 10.090 ;
        RECT 38.840 8.690 40.540 10.090 ;
        RECT 40.840 8.690 42.540 10.090 ;
        RECT 42.840 8.690 44.540 10.090 ;
        RECT 44.840 8.690 46.540 10.090 ;
        RECT 46.840 8.690 48.540 10.090 ;
        RECT 48.840 8.690 50.540 10.090 ;
        RECT 50.840 8.690 52.540 10.090 ;
        RECT 52.840 8.690 54.540 10.090 ;
        RECT 54.840 8.690 56.540 10.090 ;
        RECT 56.840 8.690 58.540 10.090 ;
        RECT 58.840 8.690 60.540 10.090 ;
        RECT 60.840 8.690 62.540 10.090 ;
        RECT 62.840 8.690 64.540 10.090 ;
        RECT 64.840 8.690 66.540 10.090 ;
        RECT 66.840 8.690 68.540 10.090 ;
        RECT 68.840 8.690 70.540 10.090 ;
        RECT 70.840 8.690 72.540 10.090 ;
        RECT 72.840 8.690 74.540 10.090 ;
        RECT 86.575 8.690 88.275 10.090 ;
        RECT 88.575 8.690 90.275 10.090 ;
        RECT 90.575 8.690 92.275 10.090 ;
        RECT 92.575 8.690 94.275 10.090 ;
        RECT 94.575 8.690 96.275 10.090 ;
        RECT 96.575 8.690 98.275 10.090 ;
        RECT 98.575 8.690 100.275 10.090 ;
        RECT 100.575 8.690 102.275 10.090 ;
        RECT 102.575 8.690 104.275 10.090 ;
        RECT 104.575 8.690 106.275 10.090 ;
        RECT 106.575 8.690 108.275 10.090 ;
        RECT 108.575 8.690 110.275 10.090 ;
        RECT 110.575 8.690 112.275 10.090 ;
        RECT 112.575 8.690 114.275 10.090 ;
        RECT 114.575 8.690 116.275 10.090 ;
        RECT 116.575 8.690 118.275 10.090 ;
        RECT 118.575 8.690 120.275 10.090 ;
        RECT 120.575 8.690 122.275 10.090 ;
        RECT 122.575 8.690 124.275 10.090 ;
        RECT 124.575 8.690 126.275 10.090 ;
        RECT 126.575 8.690 128.275 10.090 ;
        RECT 128.575 8.690 130.275 10.090 ;
        RECT 130.575 8.690 132.275 10.090 ;
        RECT 132.575 8.690 134.275 10.090 ;
        RECT 134.575 8.690 136.275 10.090 ;
        RECT 136.575 8.690 138.275 10.090 ;
        RECT 138.575 8.690 140.275 10.090 ;
        RECT 140.575 8.690 142.275 10.090 ;
        RECT 142.575 8.690 144.275 10.090 ;
        RECT 144.575 8.690 146.275 10.090 ;
        RECT 146.575 8.690 148.275 10.090 ;
        RECT 148.575 8.690 150.275 10.090 ;
        RECT 150.575 8.690 152.275 10.090 ;
        RECT 152.575 8.690 154.275 10.090 ;
        RECT 6.840 6.840 8.540 8.240 ;
        RECT 8.840 6.840 10.540 8.240 ;
        RECT 10.840 6.840 12.540 8.240 ;
        RECT 12.840 6.840 14.540 8.240 ;
        RECT 14.840 6.840 16.540 8.240 ;
        RECT 16.840 6.840 18.540 8.240 ;
        RECT 18.840 6.840 20.540 8.240 ;
        RECT 20.840 6.840 22.540 8.240 ;
        RECT 22.840 6.840 24.540 8.240 ;
        RECT 24.840 6.840 26.540 8.240 ;
        RECT 26.840 6.840 28.540 8.240 ;
        RECT 28.840 6.840 30.540 8.240 ;
        RECT 30.840 6.840 32.540 8.240 ;
        RECT 32.840 6.840 34.540 8.240 ;
        RECT 34.840 6.840 36.540 8.240 ;
        RECT 36.840 6.840 38.540 8.240 ;
        RECT 38.840 6.840 40.540 8.240 ;
        RECT 40.840 6.840 42.540 8.240 ;
        RECT 42.840 6.840 44.540 8.240 ;
        RECT 44.840 6.840 46.540 8.240 ;
        RECT 46.840 6.840 48.540 8.240 ;
        RECT 48.840 6.840 50.540 8.240 ;
        RECT 50.840 6.840 52.540 8.240 ;
        RECT 52.840 6.840 54.540 8.240 ;
        RECT 54.840 6.840 56.540 8.240 ;
        RECT 56.840 6.840 58.540 8.240 ;
        RECT 58.840 6.840 60.540 8.240 ;
        RECT 60.840 6.840 62.540 8.240 ;
        RECT 62.840 6.840 64.540 8.240 ;
        RECT 64.840 6.840 66.540 8.240 ;
        RECT 66.840 6.840 68.540 8.240 ;
        RECT 68.840 6.840 70.540 8.240 ;
        RECT 70.840 6.840 72.540 8.240 ;
        RECT 72.840 6.840 74.540 8.240 ;
        RECT 86.575 6.840 88.275 8.240 ;
        RECT 88.575 6.840 90.275 8.240 ;
        RECT 90.575 6.840 92.275 8.240 ;
        RECT 92.575 6.840 94.275 8.240 ;
        RECT 94.575 6.840 96.275 8.240 ;
        RECT 96.575 6.840 98.275 8.240 ;
        RECT 98.575 6.840 100.275 8.240 ;
        RECT 100.575 6.840 102.275 8.240 ;
        RECT 102.575 6.840 104.275 8.240 ;
        RECT 104.575 6.840 106.275 8.240 ;
        RECT 106.575 6.840 108.275 8.240 ;
        RECT 108.575 6.840 110.275 8.240 ;
        RECT 110.575 6.840 112.275 8.240 ;
        RECT 112.575 6.840 114.275 8.240 ;
        RECT 114.575 6.840 116.275 8.240 ;
        RECT 116.575 6.840 118.275 8.240 ;
        RECT 118.575 6.840 120.275 8.240 ;
        RECT 120.575 6.840 122.275 8.240 ;
        RECT 122.575 6.840 124.275 8.240 ;
        RECT 124.575 6.840 126.275 8.240 ;
        RECT 126.575 6.840 128.275 8.240 ;
        RECT 128.575 6.840 130.275 8.240 ;
        RECT 130.575 6.840 132.275 8.240 ;
        RECT 132.575 6.840 134.275 8.240 ;
        RECT 134.575 6.840 136.275 8.240 ;
        RECT 136.575 6.840 138.275 8.240 ;
        RECT 138.575 6.840 140.275 8.240 ;
        RECT 140.575 6.840 142.275 8.240 ;
        RECT 142.575 6.840 144.275 8.240 ;
        RECT 144.575 6.840 146.275 8.240 ;
        RECT 146.575 6.840 148.275 8.240 ;
        RECT 148.575 6.840 150.275 8.240 ;
        RECT 150.575 6.840 152.275 8.240 ;
        RECT 152.575 6.840 154.275 8.240 ;
        RECT 6.840 4.990 8.540 6.390 ;
        RECT 8.840 4.990 10.540 6.390 ;
        RECT 10.840 4.990 12.540 6.390 ;
        RECT 12.840 4.990 14.540 6.390 ;
        RECT 14.840 4.990 16.540 6.390 ;
        RECT 16.840 4.990 18.540 6.390 ;
        RECT 18.840 4.990 20.540 6.390 ;
        RECT 20.840 4.990 22.540 6.390 ;
        RECT 22.840 4.990 24.540 6.390 ;
        RECT 24.840 4.990 26.540 6.390 ;
        RECT 26.840 4.990 28.540 6.390 ;
        RECT 28.840 4.990 30.540 6.390 ;
        RECT 30.840 4.990 32.540 6.390 ;
        RECT 32.840 4.990 34.540 6.390 ;
        RECT 34.840 4.990 36.540 6.390 ;
        RECT 36.840 4.990 38.540 6.390 ;
        RECT 38.840 4.990 40.540 6.390 ;
        RECT 40.840 4.990 42.540 6.390 ;
        RECT 42.840 4.990 44.540 6.390 ;
        RECT 44.840 4.990 46.540 6.390 ;
        RECT 46.840 4.990 48.540 6.390 ;
        RECT 48.840 4.990 50.540 6.390 ;
        RECT 50.840 4.990 52.540 6.390 ;
        RECT 52.840 4.990 54.540 6.390 ;
        RECT 54.840 4.990 56.540 6.390 ;
        RECT 56.840 4.990 58.540 6.390 ;
        RECT 58.840 4.990 60.540 6.390 ;
        RECT 60.840 4.990 62.540 6.390 ;
        RECT 62.840 4.990 64.540 6.390 ;
        RECT 64.840 4.990 66.540 6.390 ;
        RECT 66.840 4.990 68.540 6.390 ;
        RECT 68.840 4.990 70.540 6.390 ;
        RECT 70.840 4.990 72.540 6.390 ;
        RECT 72.840 4.990 74.540 6.390 ;
        RECT 86.575 4.990 88.275 6.390 ;
        RECT 88.575 4.990 90.275 6.390 ;
        RECT 90.575 4.990 92.275 6.390 ;
        RECT 92.575 4.990 94.275 6.390 ;
        RECT 94.575 4.990 96.275 6.390 ;
        RECT 96.575 4.990 98.275 6.390 ;
        RECT 98.575 4.990 100.275 6.390 ;
        RECT 100.575 4.990 102.275 6.390 ;
        RECT 102.575 4.990 104.275 6.390 ;
        RECT 104.575 4.990 106.275 6.390 ;
        RECT 106.575 4.990 108.275 6.390 ;
        RECT 108.575 4.990 110.275 6.390 ;
        RECT 110.575 4.990 112.275 6.390 ;
        RECT 112.575 4.990 114.275 6.390 ;
        RECT 114.575 4.990 116.275 6.390 ;
        RECT 116.575 4.990 118.275 6.390 ;
        RECT 118.575 4.990 120.275 6.390 ;
        RECT 120.575 4.990 122.275 6.390 ;
        RECT 122.575 4.990 124.275 6.390 ;
        RECT 124.575 4.990 126.275 6.390 ;
        RECT 126.575 4.990 128.275 6.390 ;
        RECT 128.575 4.990 130.275 6.390 ;
        RECT 130.575 4.990 132.275 6.390 ;
        RECT 132.575 4.990 134.275 6.390 ;
        RECT 134.575 4.990 136.275 6.390 ;
        RECT 136.575 4.990 138.275 6.390 ;
        RECT 138.575 4.990 140.275 6.390 ;
        RECT 140.575 4.990 142.275 6.390 ;
        RECT 142.575 4.990 144.275 6.390 ;
        RECT 144.575 4.990 146.275 6.390 ;
        RECT 146.575 4.990 148.275 6.390 ;
        RECT 148.575 4.990 150.275 6.390 ;
        RECT 150.575 4.990 152.275 6.390 ;
        RECT 152.575 4.990 154.275 6.390 ;
        RECT 155.575 4.690 155.875 137.590 ;
        RECT 5.240 4.390 155.875 4.690 ;
        RECT 154.225 4.340 155.175 4.390 ;
        RECT 156.225 4.040 156.525 138.215 ;
        RECT 156.875 136.515 157.175 136.690 ;
        RECT 156.825 136.165 157.225 136.515 ;
        RECT 4.590 3.740 156.525 4.040 ;
        RECT 134.290 3.690 135.240 3.740 ;
        RECT 156.875 3.390 157.175 136.165 ;
        RECT 157.525 135.865 157.825 157.615 ;
        RECT 157.475 135.515 157.875 135.865 ;
        RECT 3.940 3.090 157.175 3.390 ;
        RECT 112.210 3.040 113.160 3.090 ;
        RECT 3.290 2.150 156.850 2.450 ;
        RECT 68.050 2.100 69.000 2.150 ;
        RECT 157.525 1.550 157.825 135.515 ;
        RECT 4.000 1.250 157.825 1.550 ;
        RECT 90.130 1.200 91.080 1.250 ;
      LAYER met4 ;
        RECT 3.990 224.155 4.290 224.760 ;
        RECT 7.670 224.155 7.970 224.760 ;
        RECT 11.350 224.155 11.650 224.760 ;
        RECT 15.030 224.155 15.330 224.760 ;
        RECT 18.710 224.155 19.010 224.760 ;
        RECT 22.390 224.155 22.690 224.760 ;
        RECT 26.070 224.155 26.370 224.760 ;
        RECT 29.750 224.155 30.050 224.760 ;
        RECT 33.430 224.155 33.730 224.760 ;
        RECT 37.110 224.155 37.410 224.760 ;
        RECT 40.790 224.155 41.090 224.760 ;
        RECT 44.470 224.155 44.770 224.760 ;
        RECT 48.150 224.155 48.450 224.760 ;
        RECT 51.830 224.155 52.130 224.760 ;
        RECT 55.510 224.155 55.810 224.760 ;
        RECT 59.190 224.155 59.490 224.760 ;
        RECT 3.945 223.745 4.355 224.155 ;
        RECT 7.595 223.745 8.005 224.155 ;
        RECT 11.295 223.745 11.705 224.155 ;
        RECT 14.945 223.745 15.355 224.155 ;
        RECT 18.645 223.745 19.055 224.155 ;
        RECT 22.345 223.745 22.755 224.155 ;
        RECT 25.995 223.745 26.405 224.155 ;
        RECT 29.695 223.745 30.105 224.155 ;
        RECT 33.395 223.745 33.805 224.155 ;
        RECT 37.045 223.745 37.455 224.155 ;
        RECT 40.745 223.745 41.155 224.155 ;
        RECT 44.445 223.745 44.855 224.155 ;
        RECT 48.095 223.745 48.505 224.155 ;
        RECT 51.745 223.745 52.155 224.155 ;
        RECT 55.445 223.745 55.855 224.155 ;
        RECT 59.145 223.745 59.555 224.155 ;
        RECT 66.550 223.505 66.850 224.760 ;
        RECT 66.445 223.095 66.855 223.505 ;
        RECT 70.230 222.905 70.530 224.760 ;
        RECT 70.145 222.495 70.555 222.905 ;
        RECT 73.910 222.305 74.210 224.760 ;
        RECT 73.795 222.150 74.210 222.305 ;
        RECT 73.795 221.895 74.205 222.150 ;
        RECT 77.590 221.705 77.890 224.760 ;
        RECT 77.545 221.295 77.955 221.705 ;
        RECT 81.270 221.105 81.570 224.760 ;
        RECT 81.195 220.695 81.605 221.105 ;
        RECT 84.950 220.505 85.250 224.760 ;
        RECT 84.845 220.095 85.255 220.505 ;
        RECT 88.630 219.905 88.930 224.760 ;
        RECT 140.150 223.505 140.450 224.760 ;
        RECT 140.065 223.095 140.475 223.505 ;
        RECT 143.830 222.905 144.130 224.760 ;
        RECT 143.745 222.495 144.155 222.905 ;
        RECT 147.510 222.305 147.810 224.760 ;
        RECT 147.425 221.895 147.835 222.305 ;
        RECT 151.190 221.705 151.490 224.760 ;
        RECT 151.105 221.295 151.515 221.705 ;
        RECT 154.870 221.105 155.170 224.760 ;
        RECT 154.785 220.695 155.195 221.105 ;
        RECT 158.500 220.760 160.000 224.150 ;
        RECT 88.545 219.495 88.955 219.905 ;
        RECT 29.380 216.295 30.980 218.035 ;
        RECT 32.680 216.480 34.280 218.035 ;
        RECT 29.335 215.150 31.045 216.295 ;
        RECT 2.500 213.650 31.045 215.150 ;
        RECT 29.335 205.400 31.045 213.650 ;
        RECT 32.640 215.230 34.340 216.480 ;
        RECT 32.640 213.730 158.500 215.230 ;
        RECT 31.635 206.410 31.965 206.740 ;
        RECT 2.500 203.900 31.045 205.400 ;
        RECT 29.335 195.450 31.045 203.900 ;
        RECT 31.650 197.900 31.950 206.410 ;
        RECT 31.635 197.570 31.965 197.900 ;
        RECT 2.500 193.950 31.045 195.450 ;
        RECT 29.335 184.735 31.045 193.950 ;
        RECT 32.640 191.480 34.340 213.730 ;
        RECT 105.235 207.090 105.565 207.420 ;
        RECT 51.875 201.650 52.205 201.980 ;
        RECT 51.890 197.220 52.190 201.650 ;
        RECT 51.875 196.890 52.205 197.220 ;
        RECT 105.250 195.860 105.550 207.090 ;
        RECT 105.235 195.530 105.565 195.860 ;
        RECT 32.640 189.980 158.500 191.480 ;
        RECT 32.640 185.245 34.340 189.980 ;
        RECT 142.240 185.445 145.040 185.640 ;
        RECT 29.335 184.550 31.040 184.735 ;
        RECT 2.500 183.050 31.040 184.550 ;
        RECT 32.635 183.535 34.345 185.245 ;
        RECT 142.235 184.685 145.045 185.445 ;
        RECT 142.240 184.030 145.040 184.685 ;
        RECT 29.340 182.695 31.040 183.050 ;
        RECT 29.335 180.985 31.045 182.695 ;
        RECT 29.340 172.250 31.040 180.985 ;
        RECT 2.500 170.750 31.040 172.250 ;
        RECT 29.340 159.450 31.040 170.750 ;
        RECT 32.640 165.945 34.340 183.535 ;
        RECT 125.685 180.985 127.545 182.695 ;
        RECT 142.240 182.530 158.500 184.030 ;
        RECT 81.635 177.335 81.995 177.695 ;
        RECT 79.685 173.740 80.045 173.895 ;
        RECT 79.685 173.535 80.090 173.740 ;
        RECT 32.635 164.235 34.345 165.945 ;
        RECT 32.640 160.245 34.340 164.235 ;
        RECT 32.635 159.785 34.345 160.245 ;
        RECT 2.500 157.950 31.040 159.450 ;
        RECT 29.340 154.495 31.040 157.950 ;
        RECT 29.335 152.785 31.045 154.495 ;
        RECT 29.340 152.640 31.040 152.785 ;
        RECT 32.640 146.045 34.340 159.785 ;
        RECT 32.635 139.995 34.345 146.045 ;
        RECT 48.490 140.215 48.990 140.715 ;
        RECT 32.635 138.285 36.995 139.995 ;
        RECT 48.590 131.940 48.890 140.215 ;
        RECT 79.790 131.940 80.090 173.535 ;
        RECT 48.590 131.640 80.090 131.940 ;
        RECT 79.790 127.990 80.090 131.640 ;
        RECT 71.690 127.690 80.090 127.990 ;
        RECT 81.690 131.940 81.990 177.335 ;
        RECT 125.690 154.495 127.540 180.985 ;
        RECT 142.240 167.665 145.040 182.530 ;
        RECT 142.240 166.165 158.500 167.665 ;
        RECT 142.240 165.945 145.045 166.165 ;
        RECT 142.235 164.235 145.045 165.945 ;
        RECT 125.690 152.640 129.395 154.495 ;
        RECT 127.535 152.635 129.395 152.640 ;
        RECT 112.125 140.215 112.625 140.715 ;
        RECT 112.240 131.940 112.540 140.215 ;
        RECT 81.690 131.640 112.540 131.940 ;
        RECT 81.690 127.990 81.990 131.640 ;
        RECT 81.690 127.690 89.425 127.990 ;
        RECT 7.340 127.140 8.340 127.640 ;
        RECT 7.690 126.440 7.990 127.140 ;
        RECT 9.690 126.440 9.990 126.890 ;
        RECT 11.690 126.440 11.990 126.890 ;
        RECT 13.690 126.440 13.990 126.890 ;
        RECT 15.690 126.440 15.990 126.890 ;
        RECT 17.690 126.440 17.990 126.890 ;
        RECT 19.690 126.440 19.990 126.890 ;
        RECT 21.690 126.440 21.990 126.890 ;
        RECT 23.690 126.440 23.990 126.890 ;
        RECT 25.690 126.440 25.990 126.890 ;
        RECT 27.690 126.440 27.990 126.890 ;
        RECT 29.690 126.440 29.990 126.890 ;
        RECT 31.690 126.440 31.990 126.890 ;
        RECT 33.690 126.440 33.990 126.890 ;
        RECT 35.690 126.440 35.990 126.890 ;
        RECT 37.690 126.440 37.990 126.890 ;
        RECT 39.690 126.440 39.990 126.890 ;
        RECT 41.690 126.440 41.990 126.890 ;
        RECT 43.690 126.440 43.990 126.890 ;
        RECT 45.690 126.440 45.990 126.890 ;
        RECT 47.690 126.440 47.990 126.890 ;
        RECT 49.690 126.440 49.990 126.890 ;
        RECT 51.690 126.440 51.990 126.890 ;
        RECT 53.690 126.440 53.990 126.890 ;
        RECT 55.690 126.440 55.990 126.890 ;
        RECT 57.690 126.440 57.990 126.890 ;
        RECT 59.690 126.440 59.990 126.890 ;
        RECT 61.690 126.440 61.990 126.890 ;
        RECT 63.690 126.440 63.990 126.890 ;
        RECT 65.690 126.440 65.990 126.890 ;
        RECT 67.690 126.440 67.990 126.890 ;
        RECT 69.690 126.440 69.990 126.890 ;
        RECT 71.690 126.440 71.990 127.690 ;
        RECT 73.340 126.890 74.340 127.390 ;
        RECT 86.775 126.890 87.775 127.390 ;
        RECT 73.690 126.440 73.990 126.890 ;
        RECT 87.125 126.440 87.425 126.890 ;
        RECT 89.125 126.440 89.425 127.690 ;
        RECT 152.775 127.140 153.775 127.640 ;
        RECT 91.125 126.440 91.425 126.890 ;
        RECT 93.125 126.440 93.425 126.890 ;
        RECT 95.125 126.440 95.425 126.890 ;
        RECT 97.125 126.440 97.425 126.890 ;
        RECT 99.125 126.440 99.425 126.890 ;
        RECT 101.125 126.440 101.425 126.890 ;
        RECT 103.125 126.440 103.425 126.890 ;
        RECT 105.125 126.440 105.425 126.890 ;
        RECT 107.125 126.440 107.425 126.890 ;
        RECT 109.125 126.440 109.425 126.890 ;
        RECT 111.125 126.440 111.425 126.890 ;
        RECT 113.125 126.440 113.425 126.890 ;
        RECT 115.125 126.440 115.425 126.890 ;
        RECT 117.125 126.440 117.425 126.890 ;
        RECT 119.125 126.440 119.425 126.890 ;
        RECT 121.125 126.440 121.425 126.890 ;
        RECT 123.125 126.440 123.425 126.890 ;
        RECT 125.125 126.440 125.425 126.890 ;
        RECT 127.125 126.440 127.425 126.890 ;
        RECT 129.125 126.440 129.425 126.890 ;
        RECT 131.125 126.440 131.425 126.890 ;
        RECT 133.125 126.440 133.425 126.890 ;
        RECT 135.125 126.440 135.425 126.890 ;
        RECT 137.125 126.440 137.425 126.890 ;
        RECT 139.125 126.440 139.425 126.890 ;
        RECT 141.125 126.440 141.425 126.890 ;
        RECT 143.125 126.440 143.425 126.890 ;
        RECT 145.125 126.440 145.425 126.890 ;
        RECT 147.125 126.440 147.425 126.890 ;
        RECT 149.125 126.440 149.425 126.890 ;
        RECT 151.125 126.440 151.425 126.890 ;
        RECT 153.125 126.440 153.425 127.140 ;
        RECT 7.340 125.440 8.340 126.440 ;
        RECT 9.340 126.090 10.340 126.440 ;
        RECT 11.340 126.090 12.340 126.440 ;
        RECT 13.340 126.090 14.340 126.440 ;
        RECT 15.340 126.090 16.340 126.440 ;
        RECT 17.340 126.090 18.340 126.440 ;
        RECT 19.340 126.090 20.340 126.440 ;
        RECT 21.340 126.090 22.340 126.440 ;
        RECT 23.340 126.090 24.340 126.440 ;
        RECT 25.340 126.090 26.340 126.440 ;
        RECT 27.340 126.090 28.340 126.440 ;
        RECT 29.340 126.090 30.340 126.440 ;
        RECT 31.340 126.090 32.340 126.440 ;
        RECT 33.340 126.090 34.340 126.440 ;
        RECT 35.340 126.090 36.340 126.440 ;
        RECT 37.340 126.090 38.340 126.440 ;
        RECT 39.340 126.090 40.340 126.440 ;
        RECT 41.340 126.090 42.340 126.440 ;
        RECT 43.340 126.090 44.340 126.440 ;
        RECT 45.340 126.090 46.340 126.440 ;
        RECT 47.340 126.090 48.340 126.440 ;
        RECT 49.340 126.090 50.340 126.440 ;
        RECT 51.340 126.090 52.340 126.440 ;
        RECT 53.340 126.090 54.340 126.440 ;
        RECT 55.340 126.090 56.340 126.440 ;
        RECT 57.340 126.090 58.340 126.440 ;
        RECT 59.340 126.090 60.340 126.440 ;
        RECT 61.340 126.090 62.340 126.440 ;
        RECT 63.340 126.090 64.340 126.440 ;
        RECT 65.340 126.090 66.340 126.440 ;
        RECT 67.340 126.090 68.340 126.440 ;
        RECT 69.340 126.090 70.340 126.440 ;
        RECT 71.340 126.090 72.340 126.440 ;
        RECT 9.340 125.790 72.340 126.090 ;
        RECT 9.340 125.440 10.340 125.790 ;
        RECT 11.340 125.440 12.340 125.790 ;
        RECT 13.340 125.440 14.340 125.790 ;
        RECT 15.340 125.440 16.340 125.790 ;
        RECT 17.340 125.440 18.340 125.790 ;
        RECT 19.340 125.440 20.340 125.790 ;
        RECT 21.340 125.440 22.340 125.790 ;
        RECT 23.340 125.440 24.340 125.790 ;
        RECT 25.340 125.440 26.340 125.790 ;
        RECT 27.340 125.440 28.340 125.790 ;
        RECT 29.340 125.440 30.340 125.790 ;
        RECT 31.340 125.440 32.340 125.790 ;
        RECT 33.340 125.440 34.340 125.790 ;
        RECT 35.340 125.440 36.340 125.790 ;
        RECT 37.340 125.440 38.340 125.790 ;
        RECT 39.340 125.440 40.340 125.790 ;
        RECT 41.340 125.440 42.340 125.790 ;
        RECT 43.340 125.440 44.340 125.790 ;
        RECT 45.340 125.440 46.340 125.790 ;
        RECT 47.340 125.440 48.340 125.790 ;
        RECT 49.340 125.440 50.340 125.790 ;
        RECT 51.340 125.440 52.340 125.790 ;
        RECT 53.340 125.440 54.340 125.790 ;
        RECT 55.340 125.440 56.340 125.790 ;
        RECT 57.340 125.440 58.340 125.790 ;
        RECT 59.340 125.440 60.340 125.790 ;
        RECT 61.340 125.440 62.340 125.790 ;
        RECT 63.340 125.440 64.340 125.790 ;
        RECT 65.340 125.440 66.340 125.790 ;
        RECT 67.340 125.440 68.340 125.790 ;
        RECT 69.340 125.440 70.340 125.790 ;
        RECT 71.340 125.440 72.340 125.790 ;
        RECT 73.340 125.440 74.340 126.440 ;
        RECT 86.775 125.440 87.775 126.440 ;
        RECT 88.775 126.090 89.775 126.440 ;
        RECT 90.775 126.090 91.775 126.440 ;
        RECT 92.775 126.090 93.775 126.440 ;
        RECT 94.775 126.090 95.775 126.440 ;
        RECT 96.775 126.090 97.775 126.440 ;
        RECT 98.775 126.090 99.775 126.440 ;
        RECT 100.775 126.090 101.775 126.440 ;
        RECT 102.775 126.090 103.775 126.440 ;
        RECT 104.775 126.090 105.775 126.440 ;
        RECT 106.775 126.090 107.775 126.440 ;
        RECT 108.775 126.090 109.775 126.440 ;
        RECT 110.775 126.090 111.775 126.440 ;
        RECT 112.775 126.090 113.775 126.440 ;
        RECT 114.775 126.090 115.775 126.440 ;
        RECT 116.775 126.090 117.775 126.440 ;
        RECT 118.775 126.090 119.775 126.440 ;
        RECT 120.775 126.090 121.775 126.440 ;
        RECT 122.775 126.090 123.775 126.440 ;
        RECT 124.775 126.090 125.775 126.440 ;
        RECT 126.775 126.090 127.775 126.440 ;
        RECT 128.775 126.090 129.775 126.440 ;
        RECT 130.775 126.090 131.775 126.440 ;
        RECT 132.775 126.090 133.775 126.440 ;
        RECT 134.775 126.090 135.775 126.440 ;
        RECT 136.775 126.090 137.775 126.440 ;
        RECT 138.775 126.090 139.775 126.440 ;
        RECT 140.775 126.090 141.775 126.440 ;
        RECT 142.775 126.090 143.775 126.440 ;
        RECT 144.775 126.090 145.775 126.440 ;
        RECT 146.775 126.090 147.775 126.440 ;
        RECT 148.775 126.090 149.775 126.440 ;
        RECT 150.775 126.090 151.775 126.440 ;
        RECT 88.775 125.790 151.775 126.090 ;
        RECT 88.775 125.440 89.775 125.790 ;
        RECT 90.775 125.440 91.775 125.790 ;
        RECT 92.775 125.440 93.775 125.790 ;
        RECT 94.775 125.440 95.775 125.790 ;
        RECT 96.775 125.440 97.775 125.790 ;
        RECT 98.775 125.440 99.775 125.790 ;
        RECT 100.775 125.440 101.775 125.790 ;
        RECT 102.775 125.440 103.775 125.790 ;
        RECT 104.775 125.440 105.775 125.790 ;
        RECT 106.775 125.440 107.775 125.790 ;
        RECT 108.775 125.440 109.775 125.790 ;
        RECT 110.775 125.440 111.775 125.790 ;
        RECT 112.775 125.440 113.775 125.790 ;
        RECT 114.775 125.440 115.775 125.790 ;
        RECT 116.775 125.440 117.775 125.790 ;
        RECT 118.775 125.440 119.775 125.790 ;
        RECT 120.775 125.440 121.775 125.790 ;
        RECT 122.775 125.440 123.775 125.790 ;
        RECT 124.775 125.440 125.775 125.790 ;
        RECT 126.775 125.440 127.775 125.790 ;
        RECT 128.775 125.440 129.775 125.790 ;
        RECT 130.775 125.440 131.775 125.790 ;
        RECT 132.775 125.440 133.775 125.790 ;
        RECT 134.775 125.440 135.775 125.790 ;
        RECT 136.775 125.440 137.775 125.790 ;
        RECT 138.775 125.440 139.775 125.790 ;
        RECT 140.775 125.440 141.775 125.790 ;
        RECT 142.775 125.440 143.775 125.790 ;
        RECT 144.775 125.440 145.775 125.790 ;
        RECT 146.775 125.440 147.775 125.790 ;
        RECT 148.775 125.440 149.775 125.790 ;
        RECT 150.775 125.440 151.775 125.790 ;
        RECT 152.775 125.440 153.775 126.440 ;
        RECT 7.690 124.590 7.990 125.440 ;
        RECT 9.690 124.590 9.990 125.440 ;
        RECT 11.690 124.590 11.990 125.440 ;
        RECT 13.690 124.590 13.990 125.440 ;
        RECT 15.690 124.590 15.990 125.440 ;
        RECT 17.690 124.590 17.990 125.440 ;
        RECT 19.690 124.590 19.990 125.440 ;
        RECT 21.690 124.590 21.990 125.440 ;
        RECT 23.690 124.590 23.990 125.440 ;
        RECT 25.690 124.590 25.990 125.440 ;
        RECT 27.690 124.590 27.990 125.440 ;
        RECT 29.690 124.590 29.990 125.440 ;
        RECT 31.690 124.590 31.990 125.440 ;
        RECT 33.690 124.590 33.990 125.440 ;
        RECT 35.690 124.590 35.990 125.440 ;
        RECT 37.690 124.590 37.990 125.440 ;
        RECT 39.690 124.590 39.990 125.440 ;
        RECT 41.690 124.590 41.990 125.440 ;
        RECT 43.690 124.590 43.990 125.440 ;
        RECT 45.690 124.590 45.990 125.440 ;
        RECT 47.690 124.590 47.990 125.440 ;
        RECT 49.690 124.590 49.990 125.440 ;
        RECT 51.690 124.590 51.990 125.440 ;
        RECT 53.690 124.590 53.990 125.440 ;
        RECT 55.690 124.590 55.990 125.440 ;
        RECT 57.690 124.590 57.990 125.440 ;
        RECT 59.690 124.590 59.990 125.440 ;
        RECT 61.690 124.590 61.990 125.440 ;
        RECT 63.690 124.590 63.990 125.440 ;
        RECT 65.690 124.590 65.990 125.440 ;
        RECT 67.690 124.590 67.990 125.440 ;
        RECT 69.690 124.590 69.990 125.440 ;
        RECT 71.690 124.590 71.990 125.440 ;
        RECT 73.690 124.590 73.990 125.440 ;
        RECT 87.125 124.590 87.425 125.440 ;
        RECT 89.125 124.590 89.425 125.440 ;
        RECT 91.125 124.590 91.425 125.440 ;
        RECT 93.125 124.590 93.425 125.440 ;
        RECT 95.125 124.590 95.425 125.440 ;
        RECT 97.125 124.590 97.425 125.440 ;
        RECT 99.125 124.590 99.425 125.440 ;
        RECT 101.125 124.590 101.425 125.440 ;
        RECT 103.125 124.590 103.425 125.440 ;
        RECT 105.125 124.590 105.425 125.440 ;
        RECT 107.125 124.590 107.425 125.440 ;
        RECT 109.125 124.590 109.425 125.440 ;
        RECT 111.125 124.590 111.425 125.440 ;
        RECT 113.125 124.590 113.425 125.440 ;
        RECT 115.125 124.590 115.425 125.440 ;
        RECT 117.125 124.590 117.425 125.440 ;
        RECT 119.125 124.590 119.425 125.440 ;
        RECT 121.125 124.590 121.425 125.440 ;
        RECT 123.125 124.590 123.425 125.440 ;
        RECT 125.125 124.590 125.425 125.440 ;
        RECT 127.125 124.590 127.425 125.440 ;
        RECT 129.125 124.590 129.425 125.440 ;
        RECT 131.125 124.590 131.425 125.440 ;
        RECT 133.125 124.590 133.425 125.440 ;
        RECT 135.125 124.590 135.425 125.440 ;
        RECT 137.125 124.590 137.425 125.440 ;
        RECT 139.125 124.590 139.425 125.440 ;
        RECT 141.125 124.590 141.425 125.440 ;
        RECT 143.125 124.590 143.425 125.440 ;
        RECT 145.125 124.590 145.425 125.440 ;
        RECT 147.125 124.590 147.425 125.440 ;
        RECT 149.125 124.590 149.425 125.440 ;
        RECT 151.125 124.590 151.425 125.440 ;
        RECT 153.125 124.590 153.425 125.440 ;
        RECT 7.340 123.590 8.340 124.590 ;
        RECT 9.340 123.590 10.340 124.590 ;
        RECT 11.340 123.590 12.340 124.590 ;
        RECT 13.340 123.590 14.340 124.590 ;
        RECT 15.340 123.590 16.340 124.590 ;
        RECT 17.340 123.590 18.340 124.590 ;
        RECT 19.340 123.590 20.340 124.590 ;
        RECT 21.340 123.590 22.340 124.590 ;
        RECT 23.340 123.590 24.340 124.590 ;
        RECT 25.340 123.590 26.340 124.590 ;
        RECT 27.340 123.590 28.340 124.590 ;
        RECT 29.340 123.590 30.340 124.590 ;
        RECT 31.340 123.590 32.340 124.590 ;
        RECT 33.340 123.590 34.340 124.590 ;
        RECT 35.340 123.590 36.340 124.590 ;
        RECT 37.340 123.590 38.340 124.590 ;
        RECT 39.340 123.590 40.340 124.590 ;
        RECT 41.340 123.590 42.340 124.590 ;
        RECT 43.340 123.590 44.340 124.590 ;
        RECT 45.340 123.590 46.340 124.590 ;
        RECT 47.340 123.590 48.340 124.590 ;
        RECT 49.340 123.590 50.340 124.590 ;
        RECT 51.340 123.590 52.340 124.590 ;
        RECT 53.340 123.590 54.340 124.590 ;
        RECT 55.340 123.590 56.340 124.590 ;
        RECT 57.340 123.590 58.340 124.590 ;
        RECT 59.340 123.590 60.340 124.590 ;
        RECT 61.340 123.590 62.340 124.590 ;
        RECT 63.340 123.590 64.340 124.590 ;
        RECT 65.340 123.590 66.340 124.590 ;
        RECT 67.340 123.590 68.340 124.590 ;
        RECT 69.340 123.590 70.340 124.590 ;
        RECT 71.340 123.590 72.340 124.590 ;
        RECT 73.340 123.590 74.340 124.590 ;
        RECT 86.775 123.590 87.775 124.590 ;
        RECT 88.775 123.590 89.775 124.590 ;
        RECT 90.775 123.590 91.775 124.590 ;
        RECT 92.775 123.590 93.775 124.590 ;
        RECT 94.775 123.590 95.775 124.590 ;
        RECT 96.775 123.590 97.775 124.590 ;
        RECT 98.775 123.590 99.775 124.590 ;
        RECT 100.775 123.590 101.775 124.590 ;
        RECT 102.775 123.590 103.775 124.590 ;
        RECT 104.775 123.590 105.775 124.590 ;
        RECT 106.775 123.590 107.775 124.590 ;
        RECT 108.775 123.590 109.775 124.590 ;
        RECT 110.775 123.590 111.775 124.590 ;
        RECT 112.775 123.590 113.775 124.590 ;
        RECT 114.775 123.590 115.775 124.590 ;
        RECT 116.775 123.590 117.775 124.590 ;
        RECT 118.775 123.590 119.775 124.590 ;
        RECT 120.775 123.590 121.775 124.590 ;
        RECT 122.775 123.590 123.775 124.590 ;
        RECT 124.775 123.590 125.775 124.590 ;
        RECT 126.775 123.590 127.775 124.590 ;
        RECT 128.775 123.590 129.775 124.590 ;
        RECT 130.775 123.590 131.775 124.590 ;
        RECT 132.775 123.590 133.775 124.590 ;
        RECT 134.775 123.590 135.775 124.590 ;
        RECT 136.775 123.590 137.775 124.590 ;
        RECT 138.775 123.590 139.775 124.590 ;
        RECT 140.775 123.590 141.775 124.590 ;
        RECT 142.775 123.590 143.775 124.590 ;
        RECT 144.775 123.590 145.775 124.590 ;
        RECT 146.775 123.590 147.775 124.590 ;
        RECT 148.775 123.590 149.775 124.590 ;
        RECT 150.775 123.590 151.775 124.590 ;
        RECT 152.775 123.590 153.775 124.590 ;
        RECT 7.690 122.740 7.990 123.590 ;
        RECT 9.690 122.740 9.990 123.590 ;
        RECT 11.690 122.740 11.990 123.590 ;
        RECT 13.690 122.740 13.990 123.590 ;
        RECT 15.690 122.740 15.990 123.590 ;
        RECT 17.690 122.740 17.990 123.590 ;
        RECT 19.690 122.740 19.990 123.590 ;
        RECT 21.690 122.740 21.990 123.590 ;
        RECT 23.690 122.740 23.990 123.590 ;
        RECT 25.690 122.740 25.990 123.590 ;
        RECT 27.690 122.740 27.990 123.590 ;
        RECT 29.690 122.740 29.990 123.590 ;
        RECT 31.690 122.740 31.990 123.590 ;
        RECT 33.690 122.740 33.990 123.590 ;
        RECT 35.690 122.740 35.990 123.590 ;
        RECT 37.690 122.740 37.990 123.590 ;
        RECT 39.690 122.740 39.990 123.590 ;
        RECT 41.690 122.740 41.990 123.590 ;
        RECT 43.690 122.740 43.990 123.590 ;
        RECT 45.690 122.740 45.990 123.590 ;
        RECT 47.690 122.740 47.990 123.590 ;
        RECT 49.690 122.740 49.990 123.590 ;
        RECT 51.690 122.740 51.990 123.590 ;
        RECT 53.690 122.740 53.990 123.590 ;
        RECT 55.690 122.740 55.990 123.590 ;
        RECT 57.690 122.740 57.990 123.590 ;
        RECT 59.690 122.740 59.990 123.590 ;
        RECT 61.690 122.740 61.990 123.590 ;
        RECT 63.690 122.740 63.990 123.590 ;
        RECT 65.690 122.740 65.990 123.590 ;
        RECT 67.690 122.740 67.990 123.590 ;
        RECT 69.690 122.740 69.990 123.590 ;
        RECT 71.690 122.740 71.990 123.590 ;
        RECT 73.690 122.740 73.990 123.590 ;
        RECT 87.125 122.740 87.425 123.590 ;
        RECT 89.125 122.740 89.425 123.590 ;
        RECT 91.125 122.740 91.425 123.590 ;
        RECT 93.125 122.740 93.425 123.590 ;
        RECT 95.125 122.740 95.425 123.590 ;
        RECT 97.125 122.740 97.425 123.590 ;
        RECT 99.125 122.740 99.425 123.590 ;
        RECT 101.125 122.740 101.425 123.590 ;
        RECT 103.125 122.740 103.425 123.590 ;
        RECT 105.125 122.740 105.425 123.590 ;
        RECT 107.125 122.740 107.425 123.590 ;
        RECT 109.125 122.740 109.425 123.590 ;
        RECT 111.125 122.740 111.425 123.590 ;
        RECT 113.125 122.740 113.425 123.590 ;
        RECT 115.125 122.740 115.425 123.590 ;
        RECT 117.125 122.740 117.425 123.590 ;
        RECT 119.125 122.740 119.425 123.590 ;
        RECT 121.125 122.740 121.425 123.590 ;
        RECT 123.125 122.740 123.425 123.590 ;
        RECT 125.125 122.740 125.425 123.590 ;
        RECT 127.125 122.740 127.425 123.590 ;
        RECT 129.125 122.740 129.425 123.590 ;
        RECT 131.125 122.740 131.425 123.590 ;
        RECT 133.125 122.740 133.425 123.590 ;
        RECT 135.125 122.740 135.425 123.590 ;
        RECT 137.125 122.740 137.425 123.590 ;
        RECT 139.125 122.740 139.425 123.590 ;
        RECT 141.125 122.740 141.425 123.590 ;
        RECT 143.125 122.740 143.425 123.590 ;
        RECT 145.125 122.740 145.425 123.590 ;
        RECT 147.125 122.740 147.425 123.590 ;
        RECT 149.125 122.740 149.425 123.590 ;
        RECT 151.125 122.740 151.425 123.590 ;
        RECT 153.125 122.740 153.425 123.590 ;
        RECT 7.340 121.740 8.340 122.740 ;
        RECT 9.340 121.740 10.340 122.740 ;
        RECT 11.340 121.740 12.340 122.740 ;
        RECT 13.340 121.740 14.340 122.740 ;
        RECT 15.340 121.740 16.340 122.740 ;
        RECT 17.340 121.740 18.340 122.740 ;
        RECT 19.340 121.740 20.340 122.740 ;
        RECT 21.340 121.740 22.340 122.740 ;
        RECT 23.340 121.740 24.340 122.740 ;
        RECT 25.340 121.740 26.340 122.740 ;
        RECT 27.340 121.740 28.340 122.740 ;
        RECT 29.340 121.740 30.340 122.740 ;
        RECT 31.340 121.740 32.340 122.740 ;
        RECT 33.340 121.740 34.340 122.740 ;
        RECT 35.340 121.740 36.340 122.740 ;
        RECT 37.340 121.740 38.340 122.740 ;
        RECT 39.340 121.740 40.340 122.740 ;
        RECT 41.340 121.740 42.340 122.740 ;
        RECT 43.340 121.740 44.340 122.740 ;
        RECT 45.340 121.740 46.340 122.740 ;
        RECT 47.340 121.740 48.340 122.740 ;
        RECT 49.340 121.740 50.340 122.740 ;
        RECT 51.340 121.740 52.340 122.740 ;
        RECT 53.340 121.740 54.340 122.740 ;
        RECT 55.340 121.740 56.340 122.740 ;
        RECT 57.340 121.740 58.340 122.740 ;
        RECT 59.340 121.740 60.340 122.740 ;
        RECT 61.340 121.740 62.340 122.740 ;
        RECT 63.340 121.740 64.340 122.740 ;
        RECT 65.340 121.740 66.340 122.740 ;
        RECT 67.340 121.740 68.340 122.740 ;
        RECT 69.340 121.740 70.340 122.740 ;
        RECT 71.340 121.740 72.340 122.740 ;
        RECT 73.340 121.740 74.340 122.740 ;
        RECT 86.775 121.740 87.775 122.740 ;
        RECT 88.775 121.740 89.775 122.740 ;
        RECT 90.775 121.740 91.775 122.740 ;
        RECT 92.775 121.740 93.775 122.740 ;
        RECT 94.775 121.740 95.775 122.740 ;
        RECT 96.775 121.740 97.775 122.740 ;
        RECT 98.775 121.740 99.775 122.740 ;
        RECT 100.775 121.740 101.775 122.740 ;
        RECT 102.775 121.740 103.775 122.740 ;
        RECT 104.775 121.740 105.775 122.740 ;
        RECT 106.775 121.740 107.775 122.740 ;
        RECT 108.775 121.740 109.775 122.740 ;
        RECT 110.775 121.740 111.775 122.740 ;
        RECT 112.775 121.740 113.775 122.740 ;
        RECT 114.775 121.740 115.775 122.740 ;
        RECT 116.775 121.740 117.775 122.740 ;
        RECT 118.775 121.740 119.775 122.740 ;
        RECT 120.775 121.740 121.775 122.740 ;
        RECT 122.775 121.740 123.775 122.740 ;
        RECT 124.775 121.740 125.775 122.740 ;
        RECT 126.775 121.740 127.775 122.740 ;
        RECT 128.775 121.740 129.775 122.740 ;
        RECT 130.775 121.740 131.775 122.740 ;
        RECT 132.775 121.740 133.775 122.740 ;
        RECT 134.775 121.740 135.775 122.740 ;
        RECT 136.775 121.740 137.775 122.740 ;
        RECT 138.775 121.740 139.775 122.740 ;
        RECT 140.775 121.740 141.775 122.740 ;
        RECT 142.775 121.740 143.775 122.740 ;
        RECT 144.775 121.740 145.775 122.740 ;
        RECT 146.775 121.740 147.775 122.740 ;
        RECT 148.775 121.740 149.775 122.740 ;
        RECT 150.775 121.740 151.775 122.740 ;
        RECT 152.775 121.740 153.775 122.740 ;
        RECT 7.690 120.890 7.990 121.740 ;
        RECT 9.690 120.890 9.990 121.740 ;
        RECT 11.690 120.890 11.990 121.740 ;
        RECT 13.690 120.890 13.990 121.740 ;
        RECT 15.690 120.890 15.990 121.740 ;
        RECT 17.690 120.890 17.990 121.740 ;
        RECT 19.690 120.890 19.990 121.740 ;
        RECT 21.690 120.890 21.990 121.740 ;
        RECT 23.690 120.890 23.990 121.740 ;
        RECT 25.690 120.890 25.990 121.740 ;
        RECT 27.690 120.890 27.990 121.740 ;
        RECT 29.690 120.890 29.990 121.740 ;
        RECT 31.690 120.890 31.990 121.740 ;
        RECT 33.690 120.890 33.990 121.740 ;
        RECT 35.690 120.890 35.990 121.740 ;
        RECT 37.690 120.890 37.990 121.740 ;
        RECT 39.690 120.890 39.990 121.740 ;
        RECT 41.690 120.890 41.990 121.740 ;
        RECT 43.690 120.890 43.990 121.740 ;
        RECT 45.690 120.890 45.990 121.740 ;
        RECT 47.690 120.890 47.990 121.740 ;
        RECT 49.690 120.890 49.990 121.740 ;
        RECT 51.690 120.890 51.990 121.740 ;
        RECT 53.690 120.890 53.990 121.740 ;
        RECT 55.690 120.890 55.990 121.740 ;
        RECT 57.690 120.890 57.990 121.740 ;
        RECT 59.690 120.890 59.990 121.740 ;
        RECT 61.690 120.890 61.990 121.740 ;
        RECT 63.690 120.890 63.990 121.740 ;
        RECT 65.690 120.890 65.990 121.740 ;
        RECT 67.690 120.890 67.990 121.740 ;
        RECT 69.690 120.890 69.990 121.740 ;
        RECT 71.690 120.890 71.990 121.740 ;
        RECT 73.690 120.890 73.990 121.740 ;
        RECT 87.125 120.890 87.425 121.740 ;
        RECT 89.125 120.890 89.425 121.740 ;
        RECT 91.125 120.890 91.425 121.740 ;
        RECT 93.125 120.890 93.425 121.740 ;
        RECT 95.125 120.890 95.425 121.740 ;
        RECT 97.125 120.890 97.425 121.740 ;
        RECT 99.125 120.890 99.425 121.740 ;
        RECT 101.125 120.890 101.425 121.740 ;
        RECT 103.125 120.890 103.425 121.740 ;
        RECT 105.125 120.890 105.425 121.740 ;
        RECT 107.125 120.890 107.425 121.740 ;
        RECT 109.125 120.890 109.425 121.740 ;
        RECT 111.125 120.890 111.425 121.740 ;
        RECT 113.125 120.890 113.425 121.740 ;
        RECT 115.125 120.890 115.425 121.740 ;
        RECT 117.125 120.890 117.425 121.740 ;
        RECT 119.125 120.890 119.425 121.740 ;
        RECT 121.125 120.890 121.425 121.740 ;
        RECT 123.125 120.890 123.425 121.740 ;
        RECT 125.125 120.890 125.425 121.740 ;
        RECT 127.125 120.890 127.425 121.740 ;
        RECT 129.125 120.890 129.425 121.740 ;
        RECT 131.125 120.890 131.425 121.740 ;
        RECT 133.125 120.890 133.425 121.740 ;
        RECT 135.125 120.890 135.425 121.740 ;
        RECT 137.125 120.890 137.425 121.740 ;
        RECT 139.125 120.890 139.425 121.740 ;
        RECT 141.125 120.890 141.425 121.740 ;
        RECT 143.125 120.890 143.425 121.740 ;
        RECT 145.125 120.890 145.425 121.740 ;
        RECT 147.125 120.890 147.425 121.740 ;
        RECT 149.125 120.890 149.425 121.740 ;
        RECT 151.125 120.890 151.425 121.740 ;
        RECT 153.125 120.890 153.425 121.740 ;
        RECT 7.340 119.890 8.340 120.890 ;
        RECT 9.340 119.890 10.340 120.890 ;
        RECT 11.340 119.890 12.340 120.890 ;
        RECT 13.340 119.890 14.340 120.890 ;
        RECT 15.340 119.890 16.340 120.890 ;
        RECT 17.340 119.890 18.340 120.890 ;
        RECT 19.340 119.890 20.340 120.890 ;
        RECT 21.340 119.890 22.340 120.890 ;
        RECT 23.340 119.890 24.340 120.890 ;
        RECT 25.340 119.890 26.340 120.890 ;
        RECT 27.340 119.890 28.340 120.890 ;
        RECT 29.340 119.890 30.340 120.890 ;
        RECT 31.340 119.890 32.340 120.890 ;
        RECT 33.340 119.890 34.340 120.890 ;
        RECT 35.340 119.890 36.340 120.890 ;
        RECT 37.340 119.890 38.340 120.890 ;
        RECT 39.340 119.890 40.340 120.890 ;
        RECT 41.340 119.890 42.340 120.890 ;
        RECT 43.340 119.890 44.340 120.890 ;
        RECT 45.340 119.890 46.340 120.890 ;
        RECT 47.340 119.890 48.340 120.890 ;
        RECT 49.340 119.890 50.340 120.890 ;
        RECT 51.340 119.890 52.340 120.890 ;
        RECT 53.340 119.890 54.340 120.890 ;
        RECT 55.340 119.890 56.340 120.890 ;
        RECT 57.340 119.890 58.340 120.890 ;
        RECT 59.340 119.890 60.340 120.890 ;
        RECT 61.340 119.890 62.340 120.890 ;
        RECT 63.340 119.890 64.340 120.890 ;
        RECT 65.340 119.890 66.340 120.890 ;
        RECT 67.340 119.890 68.340 120.890 ;
        RECT 69.340 119.890 70.340 120.890 ;
        RECT 71.340 119.890 72.340 120.890 ;
        RECT 73.340 119.890 74.340 120.890 ;
        RECT 86.775 119.890 87.775 120.890 ;
        RECT 88.775 119.890 89.775 120.890 ;
        RECT 90.775 119.890 91.775 120.890 ;
        RECT 92.775 119.890 93.775 120.890 ;
        RECT 94.775 119.890 95.775 120.890 ;
        RECT 96.775 119.890 97.775 120.890 ;
        RECT 98.775 119.890 99.775 120.890 ;
        RECT 100.775 119.890 101.775 120.890 ;
        RECT 102.775 119.890 103.775 120.890 ;
        RECT 104.775 119.890 105.775 120.890 ;
        RECT 106.775 119.890 107.775 120.890 ;
        RECT 108.775 119.890 109.775 120.890 ;
        RECT 110.775 119.890 111.775 120.890 ;
        RECT 112.775 119.890 113.775 120.890 ;
        RECT 114.775 119.890 115.775 120.890 ;
        RECT 116.775 119.890 117.775 120.890 ;
        RECT 118.775 119.890 119.775 120.890 ;
        RECT 120.775 119.890 121.775 120.890 ;
        RECT 122.775 119.890 123.775 120.890 ;
        RECT 124.775 119.890 125.775 120.890 ;
        RECT 126.775 119.890 127.775 120.890 ;
        RECT 128.775 119.890 129.775 120.890 ;
        RECT 130.775 119.890 131.775 120.890 ;
        RECT 132.775 119.890 133.775 120.890 ;
        RECT 134.775 119.890 135.775 120.890 ;
        RECT 136.775 119.890 137.775 120.890 ;
        RECT 138.775 119.890 139.775 120.890 ;
        RECT 140.775 119.890 141.775 120.890 ;
        RECT 142.775 119.890 143.775 120.890 ;
        RECT 144.775 119.890 145.775 120.890 ;
        RECT 146.775 119.890 147.775 120.890 ;
        RECT 148.775 119.890 149.775 120.890 ;
        RECT 150.775 119.890 151.775 120.890 ;
        RECT 152.775 119.890 153.775 120.890 ;
        RECT 7.690 119.040 7.990 119.890 ;
        RECT 9.690 119.040 9.990 119.890 ;
        RECT 11.690 119.040 11.990 119.890 ;
        RECT 13.690 119.040 13.990 119.890 ;
        RECT 15.690 119.040 15.990 119.890 ;
        RECT 17.690 119.040 17.990 119.890 ;
        RECT 19.690 119.040 19.990 119.890 ;
        RECT 21.690 119.040 21.990 119.890 ;
        RECT 23.690 119.040 23.990 119.890 ;
        RECT 25.690 119.040 25.990 119.890 ;
        RECT 27.690 119.040 27.990 119.890 ;
        RECT 29.690 119.040 29.990 119.890 ;
        RECT 31.690 119.040 31.990 119.890 ;
        RECT 33.690 119.040 33.990 119.890 ;
        RECT 35.690 119.040 35.990 119.890 ;
        RECT 37.690 119.040 37.990 119.890 ;
        RECT 39.690 119.040 39.990 119.890 ;
        RECT 41.690 119.040 41.990 119.890 ;
        RECT 43.690 119.040 43.990 119.890 ;
        RECT 45.690 119.040 45.990 119.890 ;
        RECT 47.690 119.040 47.990 119.890 ;
        RECT 49.690 119.040 49.990 119.890 ;
        RECT 51.690 119.040 51.990 119.890 ;
        RECT 53.690 119.040 53.990 119.890 ;
        RECT 55.690 119.040 55.990 119.890 ;
        RECT 57.690 119.040 57.990 119.890 ;
        RECT 59.690 119.040 59.990 119.890 ;
        RECT 61.690 119.040 61.990 119.890 ;
        RECT 63.690 119.040 63.990 119.890 ;
        RECT 65.690 119.040 65.990 119.890 ;
        RECT 67.690 119.040 67.990 119.890 ;
        RECT 69.690 119.040 69.990 119.890 ;
        RECT 71.690 119.040 71.990 119.890 ;
        RECT 73.690 119.040 73.990 119.890 ;
        RECT 87.125 119.040 87.425 119.890 ;
        RECT 89.125 119.040 89.425 119.890 ;
        RECT 91.125 119.040 91.425 119.890 ;
        RECT 93.125 119.040 93.425 119.890 ;
        RECT 95.125 119.040 95.425 119.890 ;
        RECT 97.125 119.040 97.425 119.890 ;
        RECT 99.125 119.040 99.425 119.890 ;
        RECT 101.125 119.040 101.425 119.890 ;
        RECT 103.125 119.040 103.425 119.890 ;
        RECT 105.125 119.040 105.425 119.890 ;
        RECT 107.125 119.040 107.425 119.890 ;
        RECT 109.125 119.040 109.425 119.890 ;
        RECT 111.125 119.040 111.425 119.890 ;
        RECT 113.125 119.040 113.425 119.890 ;
        RECT 115.125 119.040 115.425 119.890 ;
        RECT 117.125 119.040 117.425 119.890 ;
        RECT 119.125 119.040 119.425 119.890 ;
        RECT 121.125 119.040 121.425 119.890 ;
        RECT 123.125 119.040 123.425 119.890 ;
        RECT 125.125 119.040 125.425 119.890 ;
        RECT 127.125 119.040 127.425 119.890 ;
        RECT 129.125 119.040 129.425 119.890 ;
        RECT 131.125 119.040 131.425 119.890 ;
        RECT 133.125 119.040 133.425 119.890 ;
        RECT 135.125 119.040 135.425 119.890 ;
        RECT 137.125 119.040 137.425 119.890 ;
        RECT 139.125 119.040 139.425 119.890 ;
        RECT 141.125 119.040 141.425 119.890 ;
        RECT 143.125 119.040 143.425 119.890 ;
        RECT 145.125 119.040 145.425 119.890 ;
        RECT 147.125 119.040 147.425 119.890 ;
        RECT 149.125 119.040 149.425 119.890 ;
        RECT 151.125 119.040 151.425 119.890 ;
        RECT 153.125 119.040 153.425 119.890 ;
        RECT 7.340 118.040 8.340 119.040 ;
        RECT 9.340 118.040 10.340 119.040 ;
        RECT 11.340 118.040 12.340 119.040 ;
        RECT 13.340 118.040 14.340 119.040 ;
        RECT 15.340 118.040 16.340 119.040 ;
        RECT 17.340 118.040 18.340 119.040 ;
        RECT 19.340 118.040 20.340 119.040 ;
        RECT 21.340 118.040 22.340 119.040 ;
        RECT 23.340 118.040 24.340 119.040 ;
        RECT 25.340 118.040 26.340 119.040 ;
        RECT 27.340 118.040 28.340 119.040 ;
        RECT 29.340 118.040 30.340 119.040 ;
        RECT 31.340 118.040 32.340 119.040 ;
        RECT 33.340 118.040 34.340 119.040 ;
        RECT 35.340 118.040 36.340 119.040 ;
        RECT 37.340 118.040 38.340 119.040 ;
        RECT 39.340 118.040 40.340 119.040 ;
        RECT 41.340 118.040 42.340 119.040 ;
        RECT 43.340 118.040 44.340 119.040 ;
        RECT 45.340 118.040 46.340 119.040 ;
        RECT 47.340 118.040 48.340 119.040 ;
        RECT 49.340 118.040 50.340 119.040 ;
        RECT 51.340 118.040 52.340 119.040 ;
        RECT 53.340 118.040 54.340 119.040 ;
        RECT 55.340 118.040 56.340 119.040 ;
        RECT 57.340 118.040 58.340 119.040 ;
        RECT 59.340 118.040 60.340 119.040 ;
        RECT 61.340 118.040 62.340 119.040 ;
        RECT 63.340 118.040 64.340 119.040 ;
        RECT 65.340 118.040 66.340 119.040 ;
        RECT 67.340 118.040 68.340 119.040 ;
        RECT 69.340 118.040 70.340 119.040 ;
        RECT 71.340 118.040 72.340 119.040 ;
        RECT 73.340 118.040 74.340 119.040 ;
        RECT 86.775 118.040 87.775 119.040 ;
        RECT 88.775 118.040 89.775 119.040 ;
        RECT 90.775 118.040 91.775 119.040 ;
        RECT 92.775 118.040 93.775 119.040 ;
        RECT 94.775 118.040 95.775 119.040 ;
        RECT 96.775 118.040 97.775 119.040 ;
        RECT 98.775 118.040 99.775 119.040 ;
        RECT 100.775 118.040 101.775 119.040 ;
        RECT 102.775 118.040 103.775 119.040 ;
        RECT 104.775 118.040 105.775 119.040 ;
        RECT 106.775 118.040 107.775 119.040 ;
        RECT 108.775 118.040 109.775 119.040 ;
        RECT 110.775 118.040 111.775 119.040 ;
        RECT 112.775 118.040 113.775 119.040 ;
        RECT 114.775 118.040 115.775 119.040 ;
        RECT 116.775 118.040 117.775 119.040 ;
        RECT 118.775 118.040 119.775 119.040 ;
        RECT 120.775 118.040 121.775 119.040 ;
        RECT 122.775 118.040 123.775 119.040 ;
        RECT 124.775 118.040 125.775 119.040 ;
        RECT 126.775 118.040 127.775 119.040 ;
        RECT 128.775 118.040 129.775 119.040 ;
        RECT 130.775 118.040 131.775 119.040 ;
        RECT 132.775 118.040 133.775 119.040 ;
        RECT 134.775 118.040 135.775 119.040 ;
        RECT 136.775 118.040 137.775 119.040 ;
        RECT 138.775 118.040 139.775 119.040 ;
        RECT 140.775 118.040 141.775 119.040 ;
        RECT 142.775 118.040 143.775 119.040 ;
        RECT 144.775 118.040 145.775 119.040 ;
        RECT 146.775 118.040 147.775 119.040 ;
        RECT 148.775 118.040 149.775 119.040 ;
        RECT 150.775 118.040 151.775 119.040 ;
        RECT 152.775 118.040 153.775 119.040 ;
        RECT 7.690 117.190 7.990 118.040 ;
        RECT 9.690 117.190 9.990 118.040 ;
        RECT 11.690 117.190 11.990 118.040 ;
        RECT 13.690 117.190 13.990 118.040 ;
        RECT 15.690 117.190 15.990 118.040 ;
        RECT 17.690 117.190 17.990 118.040 ;
        RECT 19.690 117.190 19.990 118.040 ;
        RECT 21.690 117.190 21.990 118.040 ;
        RECT 23.690 117.190 23.990 118.040 ;
        RECT 25.690 117.190 25.990 118.040 ;
        RECT 27.690 117.190 27.990 118.040 ;
        RECT 29.690 117.190 29.990 118.040 ;
        RECT 31.690 117.190 31.990 118.040 ;
        RECT 33.690 117.190 33.990 118.040 ;
        RECT 35.690 117.190 35.990 118.040 ;
        RECT 37.690 117.190 37.990 118.040 ;
        RECT 39.690 117.190 39.990 118.040 ;
        RECT 41.690 117.190 41.990 118.040 ;
        RECT 43.690 117.190 43.990 118.040 ;
        RECT 45.690 117.190 45.990 118.040 ;
        RECT 47.690 117.190 47.990 118.040 ;
        RECT 49.690 117.190 49.990 118.040 ;
        RECT 51.690 117.190 51.990 118.040 ;
        RECT 53.690 117.190 53.990 118.040 ;
        RECT 55.690 117.190 55.990 118.040 ;
        RECT 57.690 117.190 57.990 118.040 ;
        RECT 59.690 117.190 59.990 118.040 ;
        RECT 61.690 117.190 61.990 118.040 ;
        RECT 63.690 117.190 63.990 118.040 ;
        RECT 65.690 117.190 65.990 118.040 ;
        RECT 67.690 117.190 67.990 118.040 ;
        RECT 69.690 117.190 69.990 118.040 ;
        RECT 71.690 117.190 71.990 118.040 ;
        RECT 73.690 117.190 73.990 118.040 ;
        RECT 87.125 117.190 87.425 118.040 ;
        RECT 89.125 117.190 89.425 118.040 ;
        RECT 91.125 117.190 91.425 118.040 ;
        RECT 93.125 117.190 93.425 118.040 ;
        RECT 95.125 117.190 95.425 118.040 ;
        RECT 97.125 117.190 97.425 118.040 ;
        RECT 99.125 117.190 99.425 118.040 ;
        RECT 101.125 117.190 101.425 118.040 ;
        RECT 103.125 117.190 103.425 118.040 ;
        RECT 105.125 117.190 105.425 118.040 ;
        RECT 107.125 117.190 107.425 118.040 ;
        RECT 109.125 117.190 109.425 118.040 ;
        RECT 111.125 117.190 111.425 118.040 ;
        RECT 113.125 117.190 113.425 118.040 ;
        RECT 115.125 117.190 115.425 118.040 ;
        RECT 117.125 117.190 117.425 118.040 ;
        RECT 119.125 117.190 119.425 118.040 ;
        RECT 121.125 117.190 121.425 118.040 ;
        RECT 123.125 117.190 123.425 118.040 ;
        RECT 125.125 117.190 125.425 118.040 ;
        RECT 127.125 117.190 127.425 118.040 ;
        RECT 129.125 117.190 129.425 118.040 ;
        RECT 131.125 117.190 131.425 118.040 ;
        RECT 133.125 117.190 133.425 118.040 ;
        RECT 135.125 117.190 135.425 118.040 ;
        RECT 137.125 117.190 137.425 118.040 ;
        RECT 139.125 117.190 139.425 118.040 ;
        RECT 141.125 117.190 141.425 118.040 ;
        RECT 143.125 117.190 143.425 118.040 ;
        RECT 145.125 117.190 145.425 118.040 ;
        RECT 147.125 117.190 147.425 118.040 ;
        RECT 149.125 117.190 149.425 118.040 ;
        RECT 151.125 117.190 151.425 118.040 ;
        RECT 153.125 117.190 153.425 118.040 ;
        RECT 7.340 116.190 8.340 117.190 ;
        RECT 9.340 116.190 10.340 117.190 ;
        RECT 11.340 116.190 12.340 117.190 ;
        RECT 13.340 116.190 14.340 117.190 ;
        RECT 15.340 116.190 16.340 117.190 ;
        RECT 17.340 116.190 18.340 117.190 ;
        RECT 19.340 116.190 20.340 117.190 ;
        RECT 21.340 116.190 22.340 117.190 ;
        RECT 23.340 116.190 24.340 117.190 ;
        RECT 25.340 116.190 26.340 117.190 ;
        RECT 27.340 116.190 28.340 117.190 ;
        RECT 29.340 116.190 30.340 117.190 ;
        RECT 31.340 116.190 32.340 117.190 ;
        RECT 33.340 116.190 34.340 117.190 ;
        RECT 35.340 116.190 36.340 117.190 ;
        RECT 37.340 116.190 38.340 117.190 ;
        RECT 39.340 116.190 40.340 117.190 ;
        RECT 41.340 116.190 42.340 117.190 ;
        RECT 43.340 116.190 44.340 117.190 ;
        RECT 45.340 116.190 46.340 117.190 ;
        RECT 47.340 116.190 48.340 117.190 ;
        RECT 49.340 116.190 50.340 117.190 ;
        RECT 51.340 116.190 52.340 117.190 ;
        RECT 53.340 116.190 54.340 117.190 ;
        RECT 55.340 116.190 56.340 117.190 ;
        RECT 57.340 116.190 58.340 117.190 ;
        RECT 59.340 116.190 60.340 117.190 ;
        RECT 61.340 116.190 62.340 117.190 ;
        RECT 63.340 116.190 64.340 117.190 ;
        RECT 65.340 116.190 66.340 117.190 ;
        RECT 67.340 116.190 68.340 117.190 ;
        RECT 69.340 116.190 70.340 117.190 ;
        RECT 71.340 116.190 72.340 117.190 ;
        RECT 73.340 116.190 74.340 117.190 ;
        RECT 86.775 116.190 87.775 117.190 ;
        RECT 88.775 116.190 89.775 117.190 ;
        RECT 90.775 116.190 91.775 117.190 ;
        RECT 92.775 116.190 93.775 117.190 ;
        RECT 94.775 116.190 95.775 117.190 ;
        RECT 96.775 116.190 97.775 117.190 ;
        RECT 98.775 116.190 99.775 117.190 ;
        RECT 100.775 116.190 101.775 117.190 ;
        RECT 102.775 116.190 103.775 117.190 ;
        RECT 104.775 116.190 105.775 117.190 ;
        RECT 106.775 116.190 107.775 117.190 ;
        RECT 108.775 116.190 109.775 117.190 ;
        RECT 110.775 116.190 111.775 117.190 ;
        RECT 112.775 116.190 113.775 117.190 ;
        RECT 114.775 116.190 115.775 117.190 ;
        RECT 116.775 116.190 117.775 117.190 ;
        RECT 118.775 116.190 119.775 117.190 ;
        RECT 120.775 116.190 121.775 117.190 ;
        RECT 122.775 116.190 123.775 117.190 ;
        RECT 124.775 116.190 125.775 117.190 ;
        RECT 126.775 116.190 127.775 117.190 ;
        RECT 128.775 116.190 129.775 117.190 ;
        RECT 130.775 116.190 131.775 117.190 ;
        RECT 132.775 116.190 133.775 117.190 ;
        RECT 134.775 116.190 135.775 117.190 ;
        RECT 136.775 116.190 137.775 117.190 ;
        RECT 138.775 116.190 139.775 117.190 ;
        RECT 140.775 116.190 141.775 117.190 ;
        RECT 142.775 116.190 143.775 117.190 ;
        RECT 144.775 116.190 145.775 117.190 ;
        RECT 146.775 116.190 147.775 117.190 ;
        RECT 148.775 116.190 149.775 117.190 ;
        RECT 150.775 116.190 151.775 117.190 ;
        RECT 152.775 116.190 153.775 117.190 ;
        RECT 7.690 115.340 7.990 116.190 ;
        RECT 9.690 115.340 9.990 116.190 ;
        RECT 11.690 115.340 11.990 116.190 ;
        RECT 13.690 115.340 13.990 116.190 ;
        RECT 15.690 115.340 15.990 116.190 ;
        RECT 17.690 115.340 17.990 116.190 ;
        RECT 19.690 115.340 19.990 116.190 ;
        RECT 21.690 115.340 21.990 116.190 ;
        RECT 23.690 115.340 23.990 116.190 ;
        RECT 25.690 115.340 25.990 116.190 ;
        RECT 27.690 115.340 27.990 116.190 ;
        RECT 29.690 115.340 29.990 116.190 ;
        RECT 31.690 115.340 31.990 116.190 ;
        RECT 33.690 115.340 33.990 116.190 ;
        RECT 35.690 115.340 35.990 116.190 ;
        RECT 37.690 115.340 37.990 116.190 ;
        RECT 39.690 115.340 39.990 116.190 ;
        RECT 41.690 115.340 41.990 116.190 ;
        RECT 43.690 115.340 43.990 116.190 ;
        RECT 45.690 115.340 45.990 116.190 ;
        RECT 47.690 115.340 47.990 116.190 ;
        RECT 49.690 115.340 49.990 116.190 ;
        RECT 51.690 115.340 51.990 116.190 ;
        RECT 53.690 115.340 53.990 116.190 ;
        RECT 55.690 115.340 55.990 116.190 ;
        RECT 57.690 115.340 57.990 116.190 ;
        RECT 59.690 115.340 59.990 116.190 ;
        RECT 61.690 115.340 61.990 116.190 ;
        RECT 63.690 115.340 63.990 116.190 ;
        RECT 65.690 115.340 65.990 116.190 ;
        RECT 67.690 115.340 67.990 116.190 ;
        RECT 69.690 115.340 69.990 116.190 ;
        RECT 71.690 115.340 71.990 116.190 ;
        RECT 73.690 115.340 73.990 116.190 ;
        RECT 87.125 115.340 87.425 116.190 ;
        RECT 89.125 115.340 89.425 116.190 ;
        RECT 91.125 115.340 91.425 116.190 ;
        RECT 93.125 115.340 93.425 116.190 ;
        RECT 95.125 115.340 95.425 116.190 ;
        RECT 97.125 115.340 97.425 116.190 ;
        RECT 99.125 115.340 99.425 116.190 ;
        RECT 101.125 115.340 101.425 116.190 ;
        RECT 103.125 115.340 103.425 116.190 ;
        RECT 105.125 115.340 105.425 116.190 ;
        RECT 107.125 115.340 107.425 116.190 ;
        RECT 109.125 115.340 109.425 116.190 ;
        RECT 111.125 115.340 111.425 116.190 ;
        RECT 113.125 115.340 113.425 116.190 ;
        RECT 115.125 115.340 115.425 116.190 ;
        RECT 117.125 115.340 117.425 116.190 ;
        RECT 119.125 115.340 119.425 116.190 ;
        RECT 121.125 115.340 121.425 116.190 ;
        RECT 123.125 115.340 123.425 116.190 ;
        RECT 125.125 115.340 125.425 116.190 ;
        RECT 127.125 115.340 127.425 116.190 ;
        RECT 129.125 115.340 129.425 116.190 ;
        RECT 131.125 115.340 131.425 116.190 ;
        RECT 133.125 115.340 133.425 116.190 ;
        RECT 135.125 115.340 135.425 116.190 ;
        RECT 137.125 115.340 137.425 116.190 ;
        RECT 139.125 115.340 139.425 116.190 ;
        RECT 141.125 115.340 141.425 116.190 ;
        RECT 143.125 115.340 143.425 116.190 ;
        RECT 145.125 115.340 145.425 116.190 ;
        RECT 147.125 115.340 147.425 116.190 ;
        RECT 149.125 115.340 149.425 116.190 ;
        RECT 151.125 115.340 151.425 116.190 ;
        RECT 153.125 115.340 153.425 116.190 ;
        RECT 7.340 114.340 8.340 115.340 ;
        RECT 9.340 114.340 10.340 115.340 ;
        RECT 11.340 114.340 12.340 115.340 ;
        RECT 13.340 114.340 14.340 115.340 ;
        RECT 15.340 114.340 16.340 115.340 ;
        RECT 17.340 114.340 18.340 115.340 ;
        RECT 19.340 114.340 20.340 115.340 ;
        RECT 21.340 114.340 22.340 115.340 ;
        RECT 23.340 114.340 24.340 115.340 ;
        RECT 25.340 114.340 26.340 115.340 ;
        RECT 27.340 114.340 28.340 115.340 ;
        RECT 29.340 114.340 30.340 115.340 ;
        RECT 31.340 114.340 32.340 115.340 ;
        RECT 33.340 114.340 34.340 115.340 ;
        RECT 35.340 114.340 36.340 115.340 ;
        RECT 37.340 114.340 38.340 115.340 ;
        RECT 39.340 114.340 40.340 115.340 ;
        RECT 41.340 114.340 42.340 115.340 ;
        RECT 43.340 114.340 44.340 115.340 ;
        RECT 45.340 114.340 46.340 115.340 ;
        RECT 47.340 114.340 48.340 115.340 ;
        RECT 49.340 114.340 50.340 115.340 ;
        RECT 51.340 114.340 52.340 115.340 ;
        RECT 53.340 114.340 54.340 115.340 ;
        RECT 55.340 114.340 56.340 115.340 ;
        RECT 57.340 114.340 58.340 115.340 ;
        RECT 59.340 114.340 60.340 115.340 ;
        RECT 61.340 114.340 62.340 115.340 ;
        RECT 63.340 114.340 64.340 115.340 ;
        RECT 65.340 114.340 66.340 115.340 ;
        RECT 67.340 114.340 68.340 115.340 ;
        RECT 69.340 114.340 70.340 115.340 ;
        RECT 71.340 114.340 72.340 115.340 ;
        RECT 73.340 114.340 74.340 115.340 ;
        RECT 86.775 114.340 87.775 115.340 ;
        RECT 88.775 114.340 89.775 115.340 ;
        RECT 90.775 114.340 91.775 115.340 ;
        RECT 92.775 114.340 93.775 115.340 ;
        RECT 94.775 114.340 95.775 115.340 ;
        RECT 96.775 114.340 97.775 115.340 ;
        RECT 98.775 114.340 99.775 115.340 ;
        RECT 100.775 114.340 101.775 115.340 ;
        RECT 102.775 114.340 103.775 115.340 ;
        RECT 104.775 114.340 105.775 115.340 ;
        RECT 106.775 114.340 107.775 115.340 ;
        RECT 108.775 114.340 109.775 115.340 ;
        RECT 110.775 114.340 111.775 115.340 ;
        RECT 112.775 114.340 113.775 115.340 ;
        RECT 114.775 114.340 115.775 115.340 ;
        RECT 116.775 114.340 117.775 115.340 ;
        RECT 118.775 114.340 119.775 115.340 ;
        RECT 120.775 114.340 121.775 115.340 ;
        RECT 122.775 114.340 123.775 115.340 ;
        RECT 124.775 114.340 125.775 115.340 ;
        RECT 126.775 114.340 127.775 115.340 ;
        RECT 128.775 114.340 129.775 115.340 ;
        RECT 130.775 114.340 131.775 115.340 ;
        RECT 132.775 114.340 133.775 115.340 ;
        RECT 134.775 114.340 135.775 115.340 ;
        RECT 136.775 114.340 137.775 115.340 ;
        RECT 138.775 114.340 139.775 115.340 ;
        RECT 140.775 114.340 141.775 115.340 ;
        RECT 142.775 114.340 143.775 115.340 ;
        RECT 144.775 114.340 145.775 115.340 ;
        RECT 146.775 114.340 147.775 115.340 ;
        RECT 148.775 114.340 149.775 115.340 ;
        RECT 150.775 114.340 151.775 115.340 ;
        RECT 152.775 114.340 153.775 115.340 ;
        RECT 7.690 113.490 7.990 114.340 ;
        RECT 9.690 113.490 9.990 114.340 ;
        RECT 11.690 113.490 11.990 114.340 ;
        RECT 13.690 113.490 13.990 114.340 ;
        RECT 15.690 113.490 15.990 114.340 ;
        RECT 17.690 113.490 17.990 114.340 ;
        RECT 19.690 113.490 19.990 114.340 ;
        RECT 21.690 113.490 21.990 114.340 ;
        RECT 23.690 113.490 23.990 114.340 ;
        RECT 25.690 113.490 25.990 114.340 ;
        RECT 27.690 113.490 27.990 114.340 ;
        RECT 29.690 113.490 29.990 114.340 ;
        RECT 31.690 113.490 31.990 114.340 ;
        RECT 33.690 113.490 33.990 114.340 ;
        RECT 35.690 113.490 35.990 114.340 ;
        RECT 37.690 113.490 37.990 114.340 ;
        RECT 39.690 113.490 39.990 114.340 ;
        RECT 41.690 113.490 41.990 114.340 ;
        RECT 43.690 113.490 43.990 114.340 ;
        RECT 45.690 113.490 45.990 114.340 ;
        RECT 47.690 113.490 47.990 114.340 ;
        RECT 49.690 113.490 49.990 114.340 ;
        RECT 51.690 113.490 51.990 114.340 ;
        RECT 53.690 113.490 53.990 114.340 ;
        RECT 55.690 113.490 55.990 114.340 ;
        RECT 57.690 113.490 57.990 114.340 ;
        RECT 59.690 113.490 59.990 114.340 ;
        RECT 61.690 113.490 61.990 114.340 ;
        RECT 63.690 113.490 63.990 114.340 ;
        RECT 65.690 113.490 65.990 114.340 ;
        RECT 67.690 113.490 67.990 114.340 ;
        RECT 69.690 113.490 69.990 114.340 ;
        RECT 71.690 113.490 71.990 114.340 ;
        RECT 73.690 113.490 73.990 114.340 ;
        RECT 87.125 113.490 87.425 114.340 ;
        RECT 89.125 113.490 89.425 114.340 ;
        RECT 91.125 113.490 91.425 114.340 ;
        RECT 93.125 113.490 93.425 114.340 ;
        RECT 95.125 113.490 95.425 114.340 ;
        RECT 97.125 113.490 97.425 114.340 ;
        RECT 99.125 113.490 99.425 114.340 ;
        RECT 101.125 113.490 101.425 114.340 ;
        RECT 103.125 113.490 103.425 114.340 ;
        RECT 105.125 113.490 105.425 114.340 ;
        RECT 107.125 113.490 107.425 114.340 ;
        RECT 109.125 113.490 109.425 114.340 ;
        RECT 111.125 113.490 111.425 114.340 ;
        RECT 113.125 113.490 113.425 114.340 ;
        RECT 115.125 113.490 115.425 114.340 ;
        RECT 117.125 113.490 117.425 114.340 ;
        RECT 119.125 113.490 119.425 114.340 ;
        RECT 121.125 113.490 121.425 114.340 ;
        RECT 123.125 113.490 123.425 114.340 ;
        RECT 125.125 113.490 125.425 114.340 ;
        RECT 127.125 113.490 127.425 114.340 ;
        RECT 129.125 113.490 129.425 114.340 ;
        RECT 131.125 113.490 131.425 114.340 ;
        RECT 133.125 113.490 133.425 114.340 ;
        RECT 135.125 113.490 135.425 114.340 ;
        RECT 137.125 113.490 137.425 114.340 ;
        RECT 139.125 113.490 139.425 114.340 ;
        RECT 141.125 113.490 141.425 114.340 ;
        RECT 143.125 113.490 143.425 114.340 ;
        RECT 145.125 113.490 145.425 114.340 ;
        RECT 147.125 113.490 147.425 114.340 ;
        RECT 149.125 113.490 149.425 114.340 ;
        RECT 151.125 113.490 151.425 114.340 ;
        RECT 153.125 113.490 153.425 114.340 ;
        RECT 7.340 112.490 8.340 113.490 ;
        RECT 9.340 112.490 10.340 113.490 ;
        RECT 11.340 112.490 12.340 113.490 ;
        RECT 13.340 112.490 14.340 113.490 ;
        RECT 15.340 112.490 16.340 113.490 ;
        RECT 17.340 112.490 18.340 113.490 ;
        RECT 19.340 112.490 20.340 113.490 ;
        RECT 21.340 112.490 22.340 113.490 ;
        RECT 23.340 112.490 24.340 113.490 ;
        RECT 25.340 112.490 26.340 113.490 ;
        RECT 27.340 112.490 28.340 113.490 ;
        RECT 29.340 112.490 30.340 113.490 ;
        RECT 31.340 112.490 32.340 113.490 ;
        RECT 33.340 112.490 34.340 113.490 ;
        RECT 35.340 112.490 36.340 113.490 ;
        RECT 37.340 112.490 38.340 113.490 ;
        RECT 39.340 112.490 40.340 113.490 ;
        RECT 41.340 112.490 42.340 113.490 ;
        RECT 43.340 112.490 44.340 113.490 ;
        RECT 45.340 112.490 46.340 113.490 ;
        RECT 47.340 112.490 48.340 113.490 ;
        RECT 49.340 112.490 50.340 113.490 ;
        RECT 51.340 112.490 52.340 113.490 ;
        RECT 53.340 112.490 54.340 113.490 ;
        RECT 55.340 112.490 56.340 113.490 ;
        RECT 57.340 112.490 58.340 113.490 ;
        RECT 59.340 112.490 60.340 113.490 ;
        RECT 61.340 112.490 62.340 113.490 ;
        RECT 63.340 112.490 64.340 113.490 ;
        RECT 65.340 112.490 66.340 113.490 ;
        RECT 67.340 112.490 68.340 113.490 ;
        RECT 69.340 112.490 70.340 113.490 ;
        RECT 71.340 112.490 72.340 113.490 ;
        RECT 73.340 112.490 74.340 113.490 ;
        RECT 86.775 112.490 87.775 113.490 ;
        RECT 88.775 112.490 89.775 113.490 ;
        RECT 90.775 112.490 91.775 113.490 ;
        RECT 92.775 112.490 93.775 113.490 ;
        RECT 94.775 112.490 95.775 113.490 ;
        RECT 96.775 112.490 97.775 113.490 ;
        RECT 98.775 112.490 99.775 113.490 ;
        RECT 100.775 112.490 101.775 113.490 ;
        RECT 102.775 112.490 103.775 113.490 ;
        RECT 104.775 112.490 105.775 113.490 ;
        RECT 106.775 112.490 107.775 113.490 ;
        RECT 108.775 112.490 109.775 113.490 ;
        RECT 110.775 112.490 111.775 113.490 ;
        RECT 112.775 112.490 113.775 113.490 ;
        RECT 114.775 112.490 115.775 113.490 ;
        RECT 116.775 112.490 117.775 113.490 ;
        RECT 118.775 112.490 119.775 113.490 ;
        RECT 120.775 112.490 121.775 113.490 ;
        RECT 122.775 112.490 123.775 113.490 ;
        RECT 124.775 112.490 125.775 113.490 ;
        RECT 126.775 112.490 127.775 113.490 ;
        RECT 128.775 112.490 129.775 113.490 ;
        RECT 130.775 112.490 131.775 113.490 ;
        RECT 132.775 112.490 133.775 113.490 ;
        RECT 134.775 112.490 135.775 113.490 ;
        RECT 136.775 112.490 137.775 113.490 ;
        RECT 138.775 112.490 139.775 113.490 ;
        RECT 140.775 112.490 141.775 113.490 ;
        RECT 142.775 112.490 143.775 113.490 ;
        RECT 144.775 112.490 145.775 113.490 ;
        RECT 146.775 112.490 147.775 113.490 ;
        RECT 148.775 112.490 149.775 113.490 ;
        RECT 150.775 112.490 151.775 113.490 ;
        RECT 152.775 112.490 153.775 113.490 ;
        RECT 7.690 111.640 7.990 112.490 ;
        RECT 9.690 111.640 9.990 112.490 ;
        RECT 11.690 111.640 11.990 112.490 ;
        RECT 13.690 111.640 13.990 112.490 ;
        RECT 15.690 111.640 15.990 112.490 ;
        RECT 17.690 111.640 17.990 112.490 ;
        RECT 19.690 111.640 19.990 112.490 ;
        RECT 21.690 111.640 21.990 112.490 ;
        RECT 23.690 111.640 23.990 112.490 ;
        RECT 25.690 111.640 25.990 112.490 ;
        RECT 27.690 111.640 27.990 112.490 ;
        RECT 29.690 111.640 29.990 112.490 ;
        RECT 31.690 111.640 31.990 112.490 ;
        RECT 33.690 111.640 33.990 112.490 ;
        RECT 35.690 111.640 35.990 112.490 ;
        RECT 37.690 111.640 37.990 112.490 ;
        RECT 39.690 111.640 39.990 112.490 ;
        RECT 41.690 111.640 41.990 112.490 ;
        RECT 43.690 111.640 43.990 112.490 ;
        RECT 45.690 111.640 45.990 112.490 ;
        RECT 47.690 111.640 47.990 112.490 ;
        RECT 49.690 111.640 49.990 112.490 ;
        RECT 51.690 111.640 51.990 112.490 ;
        RECT 53.690 111.640 53.990 112.490 ;
        RECT 55.690 111.640 55.990 112.490 ;
        RECT 57.690 111.640 57.990 112.490 ;
        RECT 59.690 111.640 59.990 112.490 ;
        RECT 61.690 111.640 61.990 112.490 ;
        RECT 63.690 111.640 63.990 112.490 ;
        RECT 65.690 111.640 65.990 112.490 ;
        RECT 67.690 111.640 67.990 112.490 ;
        RECT 69.690 111.640 69.990 112.490 ;
        RECT 71.690 111.640 71.990 112.490 ;
        RECT 73.690 111.640 73.990 112.490 ;
        RECT 87.125 111.640 87.425 112.490 ;
        RECT 89.125 111.640 89.425 112.490 ;
        RECT 91.125 111.640 91.425 112.490 ;
        RECT 93.125 111.640 93.425 112.490 ;
        RECT 95.125 111.640 95.425 112.490 ;
        RECT 97.125 111.640 97.425 112.490 ;
        RECT 99.125 111.640 99.425 112.490 ;
        RECT 101.125 111.640 101.425 112.490 ;
        RECT 103.125 111.640 103.425 112.490 ;
        RECT 105.125 111.640 105.425 112.490 ;
        RECT 107.125 111.640 107.425 112.490 ;
        RECT 109.125 111.640 109.425 112.490 ;
        RECT 111.125 111.640 111.425 112.490 ;
        RECT 113.125 111.640 113.425 112.490 ;
        RECT 115.125 111.640 115.425 112.490 ;
        RECT 117.125 111.640 117.425 112.490 ;
        RECT 119.125 111.640 119.425 112.490 ;
        RECT 121.125 111.640 121.425 112.490 ;
        RECT 123.125 111.640 123.425 112.490 ;
        RECT 125.125 111.640 125.425 112.490 ;
        RECT 127.125 111.640 127.425 112.490 ;
        RECT 129.125 111.640 129.425 112.490 ;
        RECT 131.125 111.640 131.425 112.490 ;
        RECT 133.125 111.640 133.425 112.490 ;
        RECT 135.125 111.640 135.425 112.490 ;
        RECT 137.125 111.640 137.425 112.490 ;
        RECT 139.125 111.640 139.425 112.490 ;
        RECT 141.125 111.640 141.425 112.490 ;
        RECT 143.125 111.640 143.425 112.490 ;
        RECT 145.125 111.640 145.425 112.490 ;
        RECT 147.125 111.640 147.425 112.490 ;
        RECT 149.125 111.640 149.425 112.490 ;
        RECT 151.125 111.640 151.425 112.490 ;
        RECT 153.125 111.640 153.425 112.490 ;
        RECT 7.340 110.640 8.340 111.640 ;
        RECT 9.340 110.640 10.340 111.640 ;
        RECT 11.340 110.640 12.340 111.640 ;
        RECT 13.340 110.640 14.340 111.640 ;
        RECT 15.340 110.640 16.340 111.640 ;
        RECT 17.340 110.640 18.340 111.640 ;
        RECT 19.340 110.640 20.340 111.640 ;
        RECT 21.340 110.640 22.340 111.640 ;
        RECT 23.340 110.640 24.340 111.640 ;
        RECT 25.340 110.640 26.340 111.640 ;
        RECT 27.340 110.640 28.340 111.640 ;
        RECT 29.340 110.640 30.340 111.640 ;
        RECT 31.340 110.640 32.340 111.640 ;
        RECT 33.340 110.640 34.340 111.640 ;
        RECT 35.340 110.640 36.340 111.640 ;
        RECT 37.340 110.640 38.340 111.640 ;
        RECT 39.340 110.640 40.340 111.640 ;
        RECT 41.340 110.640 42.340 111.640 ;
        RECT 43.340 110.640 44.340 111.640 ;
        RECT 45.340 110.640 46.340 111.640 ;
        RECT 47.340 110.640 48.340 111.640 ;
        RECT 49.340 110.640 50.340 111.640 ;
        RECT 51.340 110.640 52.340 111.640 ;
        RECT 53.340 110.640 54.340 111.640 ;
        RECT 55.340 110.640 56.340 111.640 ;
        RECT 57.340 110.640 58.340 111.640 ;
        RECT 59.340 110.640 60.340 111.640 ;
        RECT 61.340 110.640 62.340 111.640 ;
        RECT 63.340 110.640 64.340 111.640 ;
        RECT 65.340 110.640 66.340 111.640 ;
        RECT 67.340 110.640 68.340 111.640 ;
        RECT 69.340 110.640 70.340 111.640 ;
        RECT 71.340 110.640 72.340 111.640 ;
        RECT 73.340 110.640 74.340 111.640 ;
        RECT 86.775 110.640 87.775 111.640 ;
        RECT 88.775 110.640 89.775 111.640 ;
        RECT 90.775 110.640 91.775 111.640 ;
        RECT 92.775 110.640 93.775 111.640 ;
        RECT 94.775 110.640 95.775 111.640 ;
        RECT 96.775 110.640 97.775 111.640 ;
        RECT 98.775 110.640 99.775 111.640 ;
        RECT 100.775 110.640 101.775 111.640 ;
        RECT 102.775 110.640 103.775 111.640 ;
        RECT 104.775 110.640 105.775 111.640 ;
        RECT 106.775 110.640 107.775 111.640 ;
        RECT 108.775 110.640 109.775 111.640 ;
        RECT 110.775 110.640 111.775 111.640 ;
        RECT 112.775 110.640 113.775 111.640 ;
        RECT 114.775 110.640 115.775 111.640 ;
        RECT 116.775 110.640 117.775 111.640 ;
        RECT 118.775 110.640 119.775 111.640 ;
        RECT 120.775 110.640 121.775 111.640 ;
        RECT 122.775 110.640 123.775 111.640 ;
        RECT 124.775 110.640 125.775 111.640 ;
        RECT 126.775 110.640 127.775 111.640 ;
        RECT 128.775 110.640 129.775 111.640 ;
        RECT 130.775 110.640 131.775 111.640 ;
        RECT 132.775 110.640 133.775 111.640 ;
        RECT 134.775 110.640 135.775 111.640 ;
        RECT 136.775 110.640 137.775 111.640 ;
        RECT 138.775 110.640 139.775 111.640 ;
        RECT 140.775 110.640 141.775 111.640 ;
        RECT 142.775 110.640 143.775 111.640 ;
        RECT 144.775 110.640 145.775 111.640 ;
        RECT 146.775 110.640 147.775 111.640 ;
        RECT 148.775 110.640 149.775 111.640 ;
        RECT 150.775 110.640 151.775 111.640 ;
        RECT 152.775 110.640 153.775 111.640 ;
        RECT 7.690 109.790 7.990 110.640 ;
        RECT 9.690 109.790 9.990 110.640 ;
        RECT 11.690 109.790 11.990 110.640 ;
        RECT 13.690 109.790 13.990 110.640 ;
        RECT 15.690 109.790 15.990 110.640 ;
        RECT 17.690 109.790 17.990 110.640 ;
        RECT 19.690 109.790 19.990 110.640 ;
        RECT 21.690 109.790 21.990 110.640 ;
        RECT 23.690 109.790 23.990 110.640 ;
        RECT 25.690 109.790 25.990 110.640 ;
        RECT 27.690 109.790 27.990 110.640 ;
        RECT 29.690 109.790 29.990 110.640 ;
        RECT 31.690 109.790 31.990 110.640 ;
        RECT 33.690 109.790 33.990 110.640 ;
        RECT 35.690 109.790 35.990 110.640 ;
        RECT 37.690 109.790 37.990 110.640 ;
        RECT 39.690 109.790 39.990 110.640 ;
        RECT 41.690 109.790 41.990 110.640 ;
        RECT 43.690 109.790 43.990 110.640 ;
        RECT 45.690 109.790 45.990 110.640 ;
        RECT 47.690 109.790 47.990 110.640 ;
        RECT 49.690 109.790 49.990 110.640 ;
        RECT 51.690 109.790 51.990 110.640 ;
        RECT 53.690 109.790 53.990 110.640 ;
        RECT 55.690 109.790 55.990 110.640 ;
        RECT 57.690 109.790 57.990 110.640 ;
        RECT 59.690 109.790 59.990 110.640 ;
        RECT 61.690 109.790 61.990 110.640 ;
        RECT 63.690 109.790 63.990 110.640 ;
        RECT 65.690 109.790 65.990 110.640 ;
        RECT 67.690 109.790 67.990 110.640 ;
        RECT 69.690 109.790 69.990 110.640 ;
        RECT 71.690 109.790 71.990 110.640 ;
        RECT 73.690 109.790 73.990 110.640 ;
        RECT 87.125 109.790 87.425 110.640 ;
        RECT 89.125 109.790 89.425 110.640 ;
        RECT 91.125 109.790 91.425 110.640 ;
        RECT 93.125 109.790 93.425 110.640 ;
        RECT 95.125 109.790 95.425 110.640 ;
        RECT 97.125 109.790 97.425 110.640 ;
        RECT 99.125 109.790 99.425 110.640 ;
        RECT 101.125 109.790 101.425 110.640 ;
        RECT 103.125 109.790 103.425 110.640 ;
        RECT 105.125 109.790 105.425 110.640 ;
        RECT 107.125 109.790 107.425 110.640 ;
        RECT 109.125 109.790 109.425 110.640 ;
        RECT 111.125 109.790 111.425 110.640 ;
        RECT 113.125 109.790 113.425 110.640 ;
        RECT 115.125 109.790 115.425 110.640 ;
        RECT 117.125 109.790 117.425 110.640 ;
        RECT 119.125 109.790 119.425 110.640 ;
        RECT 121.125 109.790 121.425 110.640 ;
        RECT 123.125 109.790 123.425 110.640 ;
        RECT 125.125 109.790 125.425 110.640 ;
        RECT 127.125 109.790 127.425 110.640 ;
        RECT 129.125 109.790 129.425 110.640 ;
        RECT 131.125 109.790 131.425 110.640 ;
        RECT 133.125 109.790 133.425 110.640 ;
        RECT 135.125 109.790 135.425 110.640 ;
        RECT 137.125 109.790 137.425 110.640 ;
        RECT 139.125 109.790 139.425 110.640 ;
        RECT 141.125 109.790 141.425 110.640 ;
        RECT 143.125 109.790 143.425 110.640 ;
        RECT 145.125 109.790 145.425 110.640 ;
        RECT 147.125 109.790 147.425 110.640 ;
        RECT 149.125 109.790 149.425 110.640 ;
        RECT 151.125 109.790 151.425 110.640 ;
        RECT 153.125 109.790 153.425 110.640 ;
        RECT 7.340 108.790 8.340 109.790 ;
        RECT 9.340 108.790 10.340 109.790 ;
        RECT 11.340 108.790 12.340 109.790 ;
        RECT 13.340 108.790 14.340 109.790 ;
        RECT 15.340 108.790 16.340 109.790 ;
        RECT 17.340 108.790 18.340 109.790 ;
        RECT 19.340 108.790 20.340 109.790 ;
        RECT 21.340 108.790 22.340 109.790 ;
        RECT 23.340 108.790 24.340 109.790 ;
        RECT 25.340 108.790 26.340 109.790 ;
        RECT 27.340 108.790 28.340 109.790 ;
        RECT 29.340 108.790 30.340 109.790 ;
        RECT 31.340 108.790 32.340 109.790 ;
        RECT 33.340 108.790 34.340 109.790 ;
        RECT 35.340 108.790 36.340 109.790 ;
        RECT 37.340 108.790 38.340 109.790 ;
        RECT 39.340 108.790 40.340 109.790 ;
        RECT 41.340 108.790 42.340 109.790 ;
        RECT 43.340 108.790 44.340 109.790 ;
        RECT 45.340 108.790 46.340 109.790 ;
        RECT 47.340 108.790 48.340 109.790 ;
        RECT 49.340 108.790 50.340 109.790 ;
        RECT 51.340 108.790 52.340 109.790 ;
        RECT 53.340 108.790 54.340 109.790 ;
        RECT 55.340 108.790 56.340 109.790 ;
        RECT 57.340 108.790 58.340 109.790 ;
        RECT 59.340 108.790 60.340 109.790 ;
        RECT 61.340 108.790 62.340 109.790 ;
        RECT 63.340 108.790 64.340 109.790 ;
        RECT 65.340 108.790 66.340 109.790 ;
        RECT 67.340 108.790 68.340 109.790 ;
        RECT 69.340 108.790 70.340 109.790 ;
        RECT 71.340 108.790 72.340 109.790 ;
        RECT 73.340 108.790 74.340 109.790 ;
        RECT 86.775 108.790 87.775 109.790 ;
        RECT 88.775 108.790 89.775 109.790 ;
        RECT 90.775 108.790 91.775 109.790 ;
        RECT 92.775 108.790 93.775 109.790 ;
        RECT 94.775 108.790 95.775 109.790 ;
        RECT 96.775 108.790 97.775 109.790 ;
        RECT 98.775 108.790 99.775 109.790 ;
        RECT 100.775 108.790 101.775 109.790 ;
        RECT 102.775 108.790 103.775 109.790 ;
        RECT 104.775 108.790 105.775 109.790 ;
        RECT 106.775 108.790 107.775 109.790 ;
        RECT 108.775 108.790 109.775 109.790 ;
        RECT 110.775 108.790 111.775 109.790 ;
        RECT 112.775 108.790 113.775 109.790 ;
        RECT 114.775 108.790 115.775 109.790 ;
        RECT 116.775 108.790 117.775 109.790 ;
        RECT 118.775 108.790 119.775 109.790 ;
        RECT 120.775 108.790 121.775 109.790 ;
        RECT 122.775 108.790 123.775 109.790 ;
        RECT 124.775 108.790 125.775 109.790 ;
        RECT 126.775 108.790 127.775 109.790 ;
        RECT 128.775 108.790 129.775 109.790 ;
        RECT 130.775 108.790 131.775 109.790 ;
        RECT 132.775 108.790 133.775 109.790 ;
        RECT 134.775 108.790 135.775 109.790 ;
        RECT 136.775 108.790 137.775 109.790 ;
        RECT 138.775 108.790 139.775 109.790 ;
        RECT 140.775 108.790 141.775 109.790 ;
        RECT 142.775 108.790 143.775 109.790 ;
        RECT 144.775 108.790 145.775 109.790 ;
        RECT 146.775 108.790 147.775 109.790 ;
        RECT 148.775 108.790 149.775 109.790 ;
        RECT 150.775 108.790 151.775 109.790 ;
        RECT 152.775 108.790 153.775 109.790 ;
        RECT 7.690 107.940 7.990 108.790 ;
        RECT 9.690 107.940 9.990 108.790 ;
        RECT 11.690 107.940 11.990 108.790 ;
        RECT 13.690 107.940 13.990 108.790 ;
        RECT 15.690 107.940 15.990 108.790 ;
        RECT 17.690 107.940 17.990 108.790 ;
        RECT 19.690 107.940 19.990 108.790 ;
        RECT 21.690 107.940 21.990 108.790 ;
        RECT 23.690 107.940 23.990 108.790 ;
        RECT 25.690 107.940 25.990 108.790 ;
        RECT 27.690 107.940 27.990 108.790 ;
        RECT 29.690 107.940 29.990 108.790 ;
        RECT 31.690 107.940 31.990 108.790 ;
        RECT 33.690 107.940 33.990 108.790 ;
        RECT 35.690 107.940 35.990 108.790 ;
        RECT 37.690 107.940 37.990 108.790 ;
        RECT 39.690 107.940 39.990 108.790 ;
        RECT 41.690 107.940 41.990 108.790 ;
        RECT 43.690 107.940 43.990 108.790 ;
        RECT 45.690 107.940 45.990 108.790 ;
        RECT 47.690 107.940 47.990 108.790 ;
        RECT 49.690 107.940 49.990 108.790 ;
        RECT 51.690 107.940 51.990 108.790 ;
        RECT 53.690 107.940 53.990 108.790 ;
        RECT 55.690 107.940 55.990 108.790 ;
        RECT 57.690 107.940 57.990 108.790 ;
        RECT 59.690 107.940 59.990 108.790 ;
        RECT 61.690 107.940 61.990 108.790 ;
        RECT 63.690 107.940 63.990 108.790 ;
        RECT 65.690 107.940 65.990 108.790 ;
        RECT 67.690 107.940 67.990 108.790 ;
        RECT 69.690 107.940 69.990 108.790 ;
        RECT 71.690 107.940 71.990 108.790 ;
        RECT 73.690 107.940 73.990 108.790 ;
        RECT 87.125 107.940 87.425 108.790 ;
        RECT 89.125 107.940 89.425 108.790 ;
        RECT 91.125 107.940 91.425 108.790 ;
        RECT 93.125 107.940 93.425 108.790 ;
        RECT 95.125 107.940 95.425 108.790 ;
        RECT 97.125 107.940 97.425 108.790 ;
        RECT 99.125 107.940 99.425 108.790 ;
        RECT 101.125 107.940 101.425 108.790 ;
        RECT 103.125 107.940 103.425 108.790 ;
        RECT 105.125 107.940 105.425 108.790 ;
        RECT 107.125 107.940 107.425 108.790 ;
        RECT 109.125 107.940 109.425 108.790 ;
        RECT 111.125 107.940 111.425 108.790 ;
        RECT 113.125 107.940 113.425 108.790 ;
        RECT 115.125 107.940 115.425 108.790 ;
        RECT 117.125 107.940 117.425 108.790 ;
        RECT 119.125 107.940 119.425 108.790 ;
        RECT 121.125 107.940 121.425 108.790 ;
        RECT 123.125 107.940 123.425 108.790 ;
        RECT 125.125 107.940 125.425 108.790 ;
        RECT 127.125 107.940 127.425 108.790 ;
        RECT 129.125 107.940 129.425 108.790 ;
        RECT 131.125 107.940 131.425 108.790 ;
        RECT 133.125 107.940 133.425 108.790 ;
        RECT 135.125 107.940 135.425 108.790 ;
        RECT 137.125 107.940 137.425 108.790 ;
        RECT 139.125 107.940 139.425 108.790 ;
        RECT 141.125 107.940 141.425 108.790 ;
        RECT 143.125 107.940 143.425 108.790 ;
        RECT 145.125 107.940 145.425 108.790 ;
        RECT 147.125 107.940 147.425 108.790 ;
        RECT 149.125 107.940 149.425 108.790 ;
        RECT 151.125 107.940 151.425 108.790 ;
        RECT 153.125 107.940 153.425 108.790 ;
        RECT 7.340 106.940 8.340 107.940 ;
        RECT 9.340 106.940 10.340 107.940 ;
        RECT 11.340 106.940 12.340 107.940 ;
        RECT 13.340 106.940 14.340 107.940 ;
        RECT 15.340 106.940 16.340 107.940 ;
        RECT 17.340 106.940 18.340 107.940 ;
        RECT 19.340 106.940 20.340 107.940 ;
        RECT 21.340 106.940 22.340 107.940 ;
        RECT 23.340 106.940 24.340 107.940 ;
        RECT 25.340 106.940 26.340 107.940 ;
        RECT 27.340 106.940 28.340 107.940 ;
        RECT 29.340 106.940 30.340 107.940 ;
        RECT 31.340 106.940 32.340 107.940 ;
        RECT 33.340 106.940 34.340 107.940 ;
        RECT 35.340 106.940 36.340 107.940 ;
        RECT 37.340 106.940 38.340 107.940 ;
        RECT 39.340 106.940 40.340 107.940 ;
        RECT 41.340 106.940 42.340 107.940 ;
        RECT 43.340 106.940 44.340 107.940 ;
        RECT 45.340 106.940 46.340 107.940 ;
        RECT 47.340 106.940 48.340 107.940 ;
        RECT 49.340 106.940 50.340 107.940 ;
        RECT 51.340 106.940 52.340 107.940 ;
        RECT 53.340 106.940 54.340 107.940 ;
        RECT 55.340 106.940 56.340 107.940 ;
        RECT 57.340 106.940 58.340 107.940 ;
        RECT 59.340 106.940 60.340 107.940 ;
        RECT 61.340 106.940 62.340 107.940 ;
        RECT 63.340 106.940 64.340 107.940 ;
        RECT 65.340 106.940 66.340 107.940 ;
        RECT 67.340 106.940 68.340 107.940 ;
        RECT 69.340 106.940 70.340 107.940 ;
        RECT 71.340 106.940 72.340 107.940 ;
        RECT 73.340 106.940 74.340 107.940 ;
        RECT 86.775 106.940 87.775 107.940 ;
        RECT 88.775 106.940 89.775 107.940 ;
        RECT 90.775 106.940 91.775 107.940 ;
        RECT 92.775 106.940 93.775 107.940 ;
        RECT 94.775 106.940 95.775 107.940 ;
        RECT 96.775 106.940 97.775 107.940 ;
        RECT 98.775 106.940 99.775 107.940 ;
        RECT 100.775 106.940 101.775 107.940 ;
        RECT 102.775 106.940 103.775 107.940 ;
        RECT 104.775 106.940 105.775 107.940 ;
        RECT 106.775 106.940 107.775 107.940 ;
        RECT 108.775 106.940 109.775 107.940 ;
        RECT 110.775 106.940 111.775 107.940 ;
        RECT 112.775 106.940 113.775 107.940 ;
        RECT 114.775 106.940 115.775 107.940 ;
        RECT 116.775 106.940 117.775 107.940 ;
        RECT 118.775 106.940 119.775 107.940 ;
        RECT 120.775 106.940 121.775 107.940 ;
        RECT 122.775 106.940 123.775 107.940 ;
        RECT 124.775 106.940 125.775 107.940 ;
        RECT 126.775 106.940 127.775 107.940 ;
        RECT 128.775 106.940 129.775 107.940 ;
        RECT 130.775 106.940 131.775 107.940 ;
        RECT 132.775 106.940 133.775 107.940 ;
        RECT 134.775 106.940 135.775 107.940 ;
        RECT 136.775 106.940 137.775 107.940 ;
        RECT 138.775 106.940 139.775 107.940 ;
        RECT 140.775 106.940 141.775 107.940 ;
        RECT 142.775 106.940 143.775 107.940 ;
        RECT 144.775 106.940 145.775 107.940 ;
        RECT 146.775 106.940 147.775 107.940 ;
        RECT 148.775 106.940 149.775 107.940 ;
        RECT 150.775 106.940 151.775 107.940 ;
        RECT 152.775 106.940 153.775 107.940 ;
        RECT 7.690 106.090 7.990 106.940 ;
        RECT 9.690 106.090 9.990 106.940 ;
        RECT 11.690 106.090 11.990 106.940 ;
        RECT 13.690 106.090 13.990 106.940 ;
        RECT 15.690 106.090 15.990 106.940 ;
        RECT 17.690 106.090 17.990 106.940 ;
        RECT 19.690 106.090 19.990 106.940 ;
        RECT 21.690 106.090 21.990 106.940 ;
        RECT 23.690 106.090 23.990 106.940 ;
        RECT 25.690 106.090 25.990 106.940 ;
        RECT 27.690 106.090 27.990 106.940 ;
        RECT 29.690 106.090 29.990 106.940 ;
        RECT 31.690 106.090 31.990 106.940 ;
        RECT 33.690 106.090 33.990 106.940 ;
        RECT 35.690 106.090 35.990 106.940 ;
        RECT 37.690 106.090 37.990 106.940 ;
        RECT 39.690 106.090 39.990 106.940 ;
        RECT 41.690 106.090 41.990 106.940 ;
        RECT 43.690 106.090 43.990 106.940 ;
        RECT 45.690 106.090 45.990 106.940 ;
        RECT 47.690 106.090 47.990 106.940 ;
        RECT 49.690 106.090 49.990 106.940 ;
        RECT 51.690 106.090 51.990 106.940 ;
        RECT 53.690 106.090 53.990 106.940 ;
        RECT 55.690 106.090 55.990 106.940 ;
        RECT 57.690 106.090 57.990 106.940 ;
        RECT 59.690 106.090 59.990 106.940 ;
        RECT 61.690 106.090 61.990 106.940 ;
        RECT 63.690 106.090 63.990 106.940 ;
        RECT 65.690 106.090 65.990 106.940 ;
        RECT 67.690 106.090 67.990 106.940 ;
        RECT 69.690 106.090 69.990 106.940 ;
        RECT 71.690 106.090 71.990 106.940 ;
        RECT 73.690 106.090 73.990 106.940 ;
        RECT 87.125 106.090 87.425 106.940 ;
        RECT 89.125 106.090 89.425 106.940 ;
        RECT 91.125 106.090 91.425 106.940 ;
        RECT 93.125 106.090 93.425 106.940 ;
        RECT 95.125 106.090 95.425 106.940 ;
        RECT 97.125 106.090 97.425 106.940 ;
        RECT 99.125 106.090 99.425 106.940 ;
        RECT 101.125 106.090 101.425 106.940 ;
        RECT 103.125 106.090 103.425 106.940 ;
        RECT 105.125 106.090 105.425 106.940 ;
        RECT 107.125 106.090 107.425 106.940 ;
        RECT 109.125 106.090 109.425 106.940 ;
        RECT 111.125 106.090 111.425 106.940 ;
        RECT 113.125 106.090 113.425 106.940 ;
        RECT 115.125 106.090 115.425 106.940 ;
        RECT 117.125 106.090 117.425 106.940 ;
        RECT 119.125 106.090 119.425 106.940 ;
        RECT 121.125 106.090 121.425 106.940 ;
        RECT 123.125 106.090 123.425 106.940 ;
        RECT 125.125 106.090 125.425 106.940 ;
        RECT 127.125 106.090 127.425 106.940 ;
        RECT 129.125 106.090 129.425 106.940 ;
        RECT 131.125 106.090 131.425 106.940 ;
        RECT 133.125 106.090 133.425 106.940 ;
        RECT 135.125 106.090 135.425 106.940 ;
        RECT 137.125 106.090 137.425 106.940 ;
        RECT 139.125 106.090 139.425 106.940 ;
        RECT 141.125 106.090 141.425 106.940 ;
        RECT 143.125 106.090 143.425 106.940 ;
        RECT 145.125 106.090 145.425 106.940 ;
        RECT 147.125 106.090 147.425 106.940 ;
        RECT 149.125 106.090 149.425 106.940 ;
        RECT 151.125 106.090 151.425 106.940 ;
        RECT 153.125 106.090 153.425 106.940 ;
        RECT 7.340 105.090 8.340 106.090 ;
        RECT 9.340 105.090 10.340 106.090 ;
        RECT 11.340 105.090 12.340 106.090 ;
        RECT 13.340 105.090 14.340 106.090 ;
        RECT 15.340 105.090 16.340 106.090 ;
        RECT 17.340 105.090 18.340 106.090 ;
        RECT 19.340 105.090 20.340 106.090 ;
        RECT 21.340 105.090 22.340 106.090 ;
        RECT 23.340 105.090 24.340 106.090 ;
        RECT 25.340 105.090 26.340 106.090 ;
        RECT 27.340 105.090 28.340 106.090 ;
        RECT 29.340 105.090 30.340 106.090 ;
        RECT 31.340 105.090 32.340 106.090 ;
        RECT 33.340 105.090 34.340 106.090 ;
        RECT 35.340 105.090 36.340 106.090 ;
        RECT 37.340 105.090 38.340 106.090 ;
        RECT 39.340 105.090 40.340 106.090 ;
        RECT 41.340 105.090 42.340 106.090 ;
        RECT 43.340 105.090 44.340 106.090 ;
        RECT 45.340 105.090 46.340 106.090 ;
        RECT 47.340 105.090 48.340 106.090 ;
        RECT 49.340 105.090 50.340 106.090 ;
        RECT 51.340 105.090 52.340 106.090 ;
        RECT 53.340 105.090 54.340 106.090 ;
        RECT 55.340 105.090 56.340 106.090 ;
        RECT 57.340 105.090 58.340 106.090 ;
        RECT 59.340 105.090 60.340 106.090 ;
        RECT 61.340 105.090 62.340 106.090 ;
        RECT 63.340 105.090 64.340 106.090 ;
        RECT 65.340 105.090 66.340 106.090 ;
        RECT 67.340 105.090 68.340 106.090 ;
        RECT 69.340 105.090 70.340 106.090 ;
        RECT 71.340 105.090 72.340 106.090 ;
        RECT 73.340 105.090 74.340 106.090 ;
        RECT 86.775 105.090 87.775 106.090 ;
        RECT 88.775 105.090 89.775 106.090 ;
        RECT 90.775 105.090 91.775 106.090 ;
        RECT 92.775 105.090 93.775 106.090 ;
        RECT 94.775 105.090 95.775 106.090 ;
        RECT 96.775 105.090 97.775 106.090 ;
        RECT 98.775 105.090 99.775 106.090 ;
        RECT 100.775 105.090 101.775 106.090 ;
        RECT 102.775 105.090 103.775 106.090 ;
        RECT 104.775 105.090 105.775 106.090 ;
        RECT 106.775 105.090 107.775 106.090 ;
        RECT 108.775 105.090 109.775 106.090 ;
        RECT 110.775 105.090 111.775 106.090 ;
        RECT 112.775 105.090 113.775 106.090 ;
        RECT 114.775 105.090 115.775 106.090 ;
        RECT 116.775 105.090 117.775 106.090 ;
        RECT 118.775 105.090 119.775 106.090 ;
        RECT 120.775 105.090 121.775 106.090 ;
        RECT 122.775 105.090 123.775 106.090 ;
        RECT 124.775 105.090 125.775 106.090 ;
        RECT 126.775 105.090 127.775 106.090 ;
        RECT 128.775 105.090 129.775 106.090 ;
        RECT 130.775 105.090 131.775 106.090 ;
        RECT 132.775 105.090 133.775 106.090 ;
        RECT 134.775 105.090 135.775 106.090 ;
        RECT 136.775 105.090 137.775 106.090 ;
        RECT 138.775 105.090 139.775 106.090 ;
        RECT 140.775 105.090 141.775 106.090 ;
        RECT 142.775 105.090 143.775 106.090 ;
        RECT 144.775 105.090 145.775 106.090 ;
        RECT 146.775 105.090 147.775 106.090 ;
        RECT 148.775 105.090 149.775 106.090 ;
        RECT 150.775 105.090 151.775 106.090 ;
        RECT 152.775 105.090 153.775 106.090 ;
        RECT 7.690 104.240 7.990 105.090 ;
        RECT 9.690 104.240 9.990 105.090 ;
        RECT 11.690 104.240 11.990 105.090 ;
        RECT 13.690 104.240 13.990 105.090 ;
        RECT 15.690 104.240 15.990 105.090 ;
        RECT 17.690 104.240 17.990 105.090 ;
        RECT 19.690 104.240 19.990 105.090 ;
        RECT 21.690 104.240 21.990 105.090 ;
        RECT 23.690 104.240 23.990 105.090 ;
        RECT 25.690 104.240 25.990 105.090 ;
        RECT 27.690 104.240 27.990 105.090 ;
        RECT 29.690 104.240 29.990 105.090 ;
        RECT 31.690 104.240 31.990 105.090 ;
        RECT 33.690 104.240 33.990 105.090 ;
        RECT 35.690 104.240 35.990 105.090 ;
        RECT 37.690 104.240 37.990 105.090 ;
        RECT 39.690 104.240 39.990 105.090 ;
        RECT 41.690 104.240 41.990 105.090 ;
        RECT 43.690 104.240 43.990 105.090 ;
        RECT 45.690 104.240 45.990 105.090 ;
        RECT 47.690 104.240 47.990 105.090 ;
        RECT 49.690 104.240 49.990 105.090 ;
        RECT 51.690 104.240 51.990 105.090 ;
        RECT 53.690 104.240 53.990 105.090 ;
        RECT 55.690 104.240 55.990 105.090 ;
        RECT 57.690 104.240 57.990 105.090 ;
        RECT 59.690 104.240 59.990 105.090 ;
        RECT 61.690 104.240 61.990 105.090 ;
        RECT 63.690 104.240 63.990 105.090 ;
        RECT 65.690 104.240 65.990 105.090 ;
        RECT 67.690 104.240 67.990 105.090 ;
        RECT 69.690 104.240 69.990 105.090 ;
        RECT 71.690 104.240 71.990 105.090 ;
        RECT 73.690 104.240 73.990 105.090 ;
        RECT 87.125 104.240 87.425 105.090 ;
        RECT 89.125 104.240 89.425 105.090 ;
        RECT 91.125 104.240 91.425 105.090 ;
        RECT 93.125 104.240 93.425 105.090 ;
        RECT 95.125 104.240 95.425 105.090 ;
        RECT 97.125 104.240 97.425 105.090 ;
        RECT 99.125 104.240 99.425 105.090 ;
        RECT 101.125 104.240 101.425 105.090 ;
        RECT 103.125 104.240 103.425 105.090 ;
        RECT 105.125 104.240 105.425 105.090 ;
        RECT 107.125 104.240 107.425 105.090 ;
        RECT 109.125 104.240 109.425 105.090 ;
        RECT 111.125 104.240 111.425 105.090 ;
        RECT 113.125 104.240 113.425 105.090 ;
        RECT 115.125 104.240 115.425 105.090 ;
        RECT 117.125 104.240 117.425 105.090 ;
        RECT 119.125 104.240 119.425 105.090 ;
        RECT 121.125 104.240 121.425 105.090 ;
        RECT 123.125 104.240 123.425 105.090 ;
        RECT 125.125 104.240 125.425 105.090 ;
        RECT 127.125 104.240 127.425 105.090 ;
        RECT 129.125 104.240 129.425 105.090 ;
        RECT 131.125 104.240 131.425 105.090 ;
        RECT 133.125 104.240 133.425 105.090 ;
        RECT 135.125 104.240 135.425 105.090 ;
        RECT 137.125 104.240 137.425 105.090 ;
        RECT 139.125 104.240 139.425 105.090 ;
        RECT 141.125 104.240 141.425 105.090 ;
        RECT 143.125 104.240 143.425 105.090 ;
        RECT 145.125 104.240 145.425 105.090 ;
        RECT 147.125 104.240 147.425 105.090 ;
        RECT 149.125 104.240 149.425 105.090 ;
        RECT 151.125 104.240 151.425 105.090 ;
        RECT 153.125 104.240 153.425 105.090 ;
        RECT 7.340 103.240 8.340 104.240 ;
        RECT 9.340 103.240 10.340 104.240 ;
        RECT 11.340 103.240 12.340 104.240 ;
        RECT 13.340 103.240 14.340 104.240 ;
        RECT 15.340 103.240 16.340 104.240 ;
        RECT 17.340 103.240 18.340 104.240 ;
        RECT 19.340 103.240 20.340 104.240 ;
        RECT 21.340 103.240 22.340 104.240 ;
        RECT 23.340 103.240 24.340 104.240 ;
        RECT 25.340 103.240 26.340 104.240 ;
        RECT 27.340 103.240 28.340 104.240 ;
        RECT 29.340 103.240 30.340 104.240 ;
        RECT 31.340 103.240 32.340 104.240 ;
        RECT 33.340 103.240 34.340 104.240 ;
        RECT 35.340 103.240 36.340 104.240 ;
        RECT 37.340 103.240 38.340 104.240 ;
        RECT 39.340 103.240 40.340 104.240 ;
        RECT 41.340 103.240 42.340 104.240 ;
        RECT 43.340 103.240 44.340 104.240 ;
        RECT 45.340 103.240 46.340 104.240 ;
        RECT 47.340 103.240 48.340 104.240 ;
        RECT 49.340 103.240 50.340 104.240 ;
        RECT 51.340 103.240 52.340 104.240 ;
        RECT 53.340 103.240 54.340 104.240 ;
        RECT 55.340 103.240 56.340 104.240 ;
        RECT 57.340 103.240 58.340 104.240 ;
        RECT 59.340 103.240 60.340 104.240 ;
        RECT 61.340 103.240 62.340 104.240 ;
        RECT 63.340 103.240 64.340 104.240 ;
        RECT 65.340 103.240 66.340 104.240 ;
        RECT 67.340 103.240 68.340 104.240 ;
        RECT 69.340 103.240 70.340 104.240 ;
        RECT 71.340 103.240 72.340 104.240 ;
        RECT 73.340 103.240 74.340 104.240 ;
        RECT 86.775 103.240 87.775 104.240 ;
        RECT 88.775 103.240 89.775 104.240 ;
        RECT 90.775 103.240 91.775 104.240 ;
        RECT 92.775 103.240 93.775 104.240 ;
        RECT 94.775 103.240 95.775 104.240 ;
        RECT 96.775 103.240 97.775 104.240 ;
        RECT 98.775 103.240 99.775 104.240 ;
        RECT 100.775 103.240 101.775 104.240 ;
        RECT 102.775 103.240 103.775 104.240 ;
        RECT 104.775 103.240 105.775 104.240 ;
        RECT 106.775 103.240 107.775 104.240 ;
        RECT 108.775 103.240 109.775 104.240 ;
        RECT 110.775 103.240 111.775 104.240 ;
        RECT 112.775 103.240 113.775 104.240 ;
        RECT 114.775 103.240 115.775 104.240 ;
        RECT 116.775 103.240 117.775 104.240 ;
        RECT 118.775 103.240 119.775 104.240 ;
        RECT 120.775 103.240 121.775 104.240 ;
        RECT 122.775 103.240 123.775 104.240 ;
        RECT 124.775 103.240 125.775 104.240 ;
        RECT 126.775 103.240 127.775 104.240 ;
        RECT 128.775 103.240 129.775 104.240 ;
        RECT 130.775 103.240 131.775 104.240 ;
        RECT 132.775 103.240 133.775 104.240 ;
        RECT 134.775 103.240 135.775 104.240 ;
        RECT 136.775 103.240 137.775 104.240 ;
        RECT 138.775 103.240 139.775 104.240 ;
        RECT 140.775 103.240 141.775 104.240 ;
        RECT 142.775 103.240 143.775 104.240 ;
        RECT 144.775 103.240 145.775 104.240 ;
        RECT 146.775 103.240 147.775 104.240 ;
        RECT 148.775 103.240 149.775 104.240 ;
        RECT 150.775 103.240 151.775 104.240 ;
        RECT 152.775 103.240 153.775 104.240 ;
        RECT 7.690 102.390 7.990 103.240 ;
        RECT 9.690 102.390 9.990 103.240 ;
        RECT 11.690 102.390 11.990 103.240 ;
        RECT 13.690 102.390 13.990 103.240 ;
        RECT 15.690 102.390 15.990 103.240 ;
        RECT 17.690 102.390 17.990 103.240 ;
        RECT 19.690 102.390 19.990 103.240 ;
        RECT 21.690 102.390 21.990 103.240 ;
        RECT 23.690 102.390 23.990 103.240 ;
        RECT 25.690 102.390 25.990 103.240 ;
        RECT 27.690 102.390 27.990 103.240 ;
        RECT 29.690 102.390 29.990 103.240 ;
        RECT 31.690 102.390 31.990 103.240 ;
        RECT 33.690 102.390 33.990 103.240 ;
        RECT 35.690 102.390 35.990 103.240 ;
        RECT 37.690 102.390 37.990 103.240 ;
        RECT 39.690 102.390 39.990 103.240 ;
        RECT 41.690 102.390 41.990 103.240 ;
        RECT 43.690 102.390 43.990 103.240 ;
        RECT 45.690 102.390 45.990 103.240 ;
        RECT 47.690 102.390 47.990 103.240 ;
        RECT 49.690 102.390 49.990 103.240 ;
        RECT 51.690 102.390 51.990 103.240 ;
        RECT 53.690 102.390 53.990 103.240 ;
        RECT 55.690 102.390 55.990 103.240 ;
        RECT 57.690 102.390 57.990 103.240 ;
        RECT 59.690 102.390 59.990 103.240 ;
        RECT 61.690 102.390 61.990 103.240 ;
        RECT 63.690 102.390 63.990 103.240 ;
        RECT 65.690 102.390 65.990 103.240 ;
        RECT 67.690 102.390 67.990 103.240 ;
        RECT 69.690 102.390 69.990 103.240 ;
        RECT 71.690 102.390 71.990 103.240 ;
        RECT 73.690 102.390 73.990 103.240 ;
        RECT 87.125 102.390 87.425 103.240 ;
        RECT 89.125 102.390 89.425 103.240 ;
        RECT 91.125 102.390 91.425 103.240 ;
        RECT 93.125 102.390 93.425 103.240 ;
        RECT 95.125 102.390 95.425 103.240 ;
        RECT 97.125 102.390 97.425 103.240 ;
        RECT 99.125 102.390 99.425 103.240 ;
        RECT 101.125 102.390 101.425 103.240 ;
        RECT 103.125 102.390 103.425 103.240 ;
        RECT 105.125 102.390 105.425 103.240 ;
        RECT 107.125 102.390 107.425 103.240 ;
        RECT 109.125 102.390 109.425 103.240 ;
        RECT 111.125 102.390 111.425 103.240 ;
        RECT 113.125 102.390 113.425 103.240 ;
        RECT 115.125 102.390 115.425 103.240 ;
        RECT 117.125 102.390 117.425 103.240 ;
        RECT 119.125 102.390 119.425 103.240 ;
        RECT 121.125 102.390 121.425 103.240 ;
        RECT 123.125 102.390 123.425 103.240 ;
        RECT 125.125 102.390 125.425 103.240 ;
        RECT 127.125 102.390 127.425 103.240 ;
        RECT 129.125 102.390 129.425 103.240 ;
        RECT 131.125 102.390 131.425 103.240 ;
        RECT 133.125 102.390 133.425 103.240 ;
        RECT 135.125 102.390 135.425 103.240 ;
        RECT 137.125 102.390 137.425 103.240 ;
        RECT 139.125 102.390 139.425 103.240 ;
        RECT 141.125 102.390 141.425 103.240 ;
        RECT 143.125 102.390 143.425 103.240 ;
        RECT 145.125 102.390 145.425 103.240 ;
        RECT 147.125 102.390 147.425 103.240 ;
        RECT 149.125 102.390 149.425 103.240 ;
        RECT 151.125 102.390 151.425 103.240 ;
        RECT 153.125 102.390 153.425 103.240 ;
        RECT 7.340 101.390 8.340 102.390 ;
        RECT 9.340 101.390 10.340 102.390 ;
        RECT 11.340 101.390 12.340 102.390 ;
        RECT 13.340 101.390 14.340 102.390 ;
        RECT 15.340 101.390 16.340 102.390 ;
        RECT 17.340 101.390 18.340 102.390 ;
        RECT 19.340 101.390 20.340 102.390 ;
        RECT 21.340 101.390 22.340 102.390 ;
        RECT 23.340 101.390 24.340 102.390 ;
        RECT 25.340 101.390 26.340 102.390 ;
        RECT 27.340 101.390 28.340 102.390 ;
        RECT 29.340 101.390 30.340 102.390 ;
        RECT 31.340 101.390 32.340 102.390 ;
        RECT 33.340 101.390 34.340 102.390 ;
        RECT 35.340 101.390 36.340 102.390 ;
        RECT 37.340 101.390 38.340 102.390 ;
        RECT 39.340 101.390 40.340 102.390 ;
        RECT 41.340 101.390 42.340 102.390 ;
        RECT 43.340 101.390 44.340 102.390 ;
        RECT 45.340 101.390 46.340 102.390 ;
        RECT 47.340 101.390 48.340 102.390 ;
        RECT 49.340 101.390 50.340 102.390 ;
        RECT 51.340 101.390 52.340 102.390 ;
        RECT 53.340 101.390 54.340 102.390 ;
        RECT 55.340 101.390 56.340 102.390 ;
        RECT 57.340 101.390 58.340 102.390 ;
        RECT 59.340 101.390 60.340 102.390 ;
        RECT 61.340 101.390 62.340 102.390 ;
        RECT 63.340 101.390 64.340 102.390 ;
        RECT 65.340 101.390 66.340 102.390 ;
        RECT 67.340 101.390 68.340 102.390 ;
        RECT 69.340 101.390 70.340 102.390 ;
        RECT 71.340 101.390 72.340 102.390 ;
        RECT 73.340 101.390 74.340 102.390 ;
        RECT 86.775 101.390 87.775 102.390 ;
        RECT 88.775 101.390 89.775 102.390 ;
        RECT 90.775 101.390 91.775 102.390 ;
        RECT 92.775 101.390 93.775 102.390 ;
        RECT 94.775 101.390 95.775 102.390 ;
        RECT 96.775 101.390 97.775 102.390 ;
        RECT 98.775 101.390 99.775 102.390 ;
        RECT 100.775 101.390 101.775 102.390 ;
        RECT 102.775 101.390 103.775 102.390 ;
        RECT 104.775 101.390 105.775 102.390 ;
        RECT 106.775 101.390 107.775 102.390 ;
        RECT 108.775 101.390 109.775 102.390 ;
        RECT 110.775 101.390 111.775 102.390 ;
        RECT 112.775 101.390 113.775 102.390 ;
        RECT 114.775 101.390 115.775 102.390 ;
        RECT 116.775 101.390 117.775 102.390 ;
        RECT 118.775 101.390 119.775 102.390 ;
        RECT 120.775 101.390 121.775 102.390 ;
        RECT 122.775 101.390 123.775 102.390 ;
        RECT 124.775 101.390 125.775 102.390 ;
        RECT 126.775 101.390 127.775 102.390 ;
        RECT 128.775 101.390 129.775 102.390 ;
        RECT 130.775 101.390 131.775 102.390 ;
        RECT 132.775 101.390 133.775 102.390 ;
        RECT 134.775 101.390 135.775 102.390 ;
        RECT 136.775 101.390 137.775 102.390 ;
        RECT 138.775 101.390 139.775 102.390 ;
        RECT 140.775 101.390 141.775 102.390 ;
        RECT 142.775 101.390 143.775 102.390 ;
        RECT 144.775 101.390 145.775 102.390 ;
        RECT 146.775 101.390 147.775 102.390 ;
        RECT 148.775 101.390 149.775 102.390 ;
        RECT 150.775 101.390 151.775 102.390 ;
        RECT 152.775 101.390 153.775 102.390 ;
        RECT 7.690 100.540 7.990 101.390 ;
        RECT 9.690 100.540 9.990 101.390 ;
        RECT 11.690 100.540 11.990 101.390 ;
        RECT 13.690 100.540 13.990 101.390 ;
        RECT 15.690 100.540 15.990 101.390 ;
        RECT 17.690 100.540 17.990 101.390 ;
        RECT 19.690 100.540 19.990 101.390 ;
        RECT 21.690 100.540 21.990 101.390 ;
        RECT 23.690 100.540 23.990 101.390 ;
        RECT 25.690 100.540 25.990 101.390 ;
        RECT 27.690 100.540 27.990 101.390 ;
        RECT 29.690 100.540 29.990 101.390 ;
        RECT 31.690 100.540 31.990 101.390 ;
        RECT 33.690 100.540 33.990 101.390 ;
        RECT 35.690 100.540 35.990 101.390 ;
        RECT 37.690 100.540 37.990 101.390 ;
        RECT 39.690 100.540 39.990 101.390 ;
        RECT 41.690 100.540 41.990 101.390 ;
        RECT 43.690 100.540 43.990 101.390 ;
        RECT 45.690 100.540 45.990 101.390 ;
        RECT 47.690 100.540 47.990 101.390 ;
        RECT 49.690 100.540 49.990 101.390 ;
        RECT 51.690 100.540 51.990 101.390 ;
        RECT 53.690 100.540 53.990 101.390 ;
        RECT 55.690 100.540 55.990 101.390 ;
        RECT 57.690 100.540 57.990 101.390 ;
        RECT 59.690 100.540 59.990 101.390 ;
        RECT 61.690 100.540 61.990 101.390 ;
        RECT 63.690 100.540 63.990 101.390 ;
        RECT 65.690 100.540 65.990 101.390 ;
        RECT 67.690 100.540 67.990 101.390 ;
        RECT 69.690 100.540 69.990 101.390 ;
        RECT 71.690 100.540 71.990 101.390 ;
        RECT 73.690 100.540 73.990 101.390 ;
        RECT 87.125 100.540 87.425 101.390 ;
        RECT 89.125 100.540 89.425 101.390 ;
        RECT 91.125 100.540 91.425 101.390 ;
        RECT 93.125 100.540 93.425 101.390 ;
        RECT 95.125 100.540 95.425 101.390 ;
        RECT 97.125 100.540 97.425 101.390 ;
        RECT 99.125 100.540 99.425 101.390 ;
        RECT 101.125 100.540 101.425 101.390 ;
        RECT 103.125 100.540 103.425 101.390 ;
        RECT 105.125 100.540 105.425 101.390 ;
        RECT 107.125 100.540 107.425 101.390 ;
        RECT 109.125 100.540 109.425 101.390 ;
        RECT 111.125 100.540 111.425 101.390 ;
        RECT 113.125 100.540 113.425 101.390 ;
        RECT 115.125 100.540 115.425 101.390 ;
        RECT 117.125 100.540 117.425 101.390 ;
        RECT 119.125 100.540 119.425 101.390 ;
        RECT 121.125 100.540 121.425 101.390 ;
        RECT 123.125 100.540 123.425 101.390 ;
        RECT 125.125 100.540 125.425 101.390 ;
        RECT 127.125 100.540 127.425 101.390 ;
        RECT 129.125 100.540 129.425 101.390 ;
        RECT 131.125 100.540 131.425 101.390 ;
        RECT 133.125 100.540 133.425 101.390 ;
        RECT 135.125 100.540 135.425 101.390 ;
        RECT 137.125 100.540 137.425 101.390 ;
        RECT 139.125 100.540 139.425 101.390 ;
        RECT 141.125 100.540 141.425 101.390 ;
        RECT 143.125 100.540 143.425 101.390 ;
        RECT 145.125 100.540 145.425 101.390 ;
        RECT 147.125 100.540 147.425 101.390 ;
        RECT 149.125 100.540 149.425 101.390 ;
        RECT 151.125 100.540 151.425 101.390 ;
        RECT 153.125 100.540 153.425 101.390 ;
        RECT 7.340 99.540 8.340 100.540 ;
        RECT 9.340 99.540 10.340 100.540 ;
        RECT 11.340 99.540 12.340 100.540 ;
        RECT 13.340 99.540 14.340 100.540 ;
        RECT 15.340 99.540 16.340 100.540 ;
        RECT 17.340 99.540 18.340 100.540 ;
        RECT 19.340 99.540 20.340 100.540 ;
        RECT 21.340 99.540 22.340 100.540 ;
        RECT 23.340 99.540 24.340 100.540 ;
        RECT 25.340 99.540 26.340 100.540 ;
        RECT 27.340 99.540 28.340 100.540 ;
        RECT 29.340 99.540 30.340 100.540 ;
        RECT 31.340 99.540 32.340 100.540 ;
        RECT 33.340 99.540 34.340 100.540 ;
        RECT 35.340 99.540 36.340 100.540 ;
        RECT 37.340 99.540 38.340 100.540 ;
        RECT 39.340 99.540 40.340 100.540 ;
        RECT 41.340 99.540 42.340 100.540 ;
        RECT 43.340 99.540 44.340 100.540 ;
        RECT 45.340 99.540 46.340 100.540 ;
        RECT 47.340 99.540 48.340 100.540 ;
        RECT 49.340 99.540 50.340 100.540 ;
        RECT 51.340 99.540 52.340 100.540 ;
        RECT 53.340 99.540 54.340 100.540 ;
        RECT 55.340 99.540 56.340 100.540 ;
        RECT 57.340 99.540 58.340 100.540 ;
        RECT 59.340 99.540 60.340 100.540 ;
        RECT 61.340 99.540 62.340 100.540 ;
        RECT 63.340 99.540 64.340 100.540 ;
        RECT 65.340 99.540 66.340 100.540 ;
        RECT 67.340 99.540 68.340 100.540 ;
        RECT 69.340 99.540 70.340 100.540 ;
        RECT 71.340 99.540 72.340 100.540 ;
        RECT 73.340 99.540 74.340 100.540 ;
        RECT 86.775 99.540 87.775 100.540 ;
        RECT 88.775 99.540 89.775 100.540 ;
        RECT 90.775 99.540 91.775 100.540 ;
        RECT 92.775 99.540 93.775 100.540 ;
        RECT 94.775 99.540 95.775 100.540 ;
        RECT 96.775 99.540 97.775 100.540 ;
        RECT 98.775 99.540 99.775 100.540 ;
        RECT 100.775 99.540 101.775 100.540 ;
        RECT 102.775 99.540 103.775 100.540 ;
        RECT 104.775 99.540 105.775 100.540 ;
        RECT 106.775 99.540 107.775 100.540 ;
        RECT 108.775 99.540 109.775 100.540 ;
        RECT 110.775 99.540 111.775 100.540 ;
        RECT 112.775 99.540 113.775 100.540 ;
        RECT 114.775 99.540 115.775 100.540 ;
        RECT 116.775 99.540 117.775 100.540 ;
        RECT 118.775 99.540 119.775 100.540 ;
        RECT 120.775 99.540 121.775 100.540 ;
        RECT 122.775 99.540 123.775 100.540 ;
        RECT 124.775 99.540 125.775 100.540 ;
        RECT 126.775 99.540 127.775 100.540 ;
        RECT 128.775 99.540 129.775 100.540 ;
        RECT 130.775 99.540 131.775 100.540 ;
        RECT 132.775 99.540 133.775 100.540 ;
        RECT 134.775 99.540 135.775 100.540 ;
        RECT 136.775 99.540 137.775 100.540 ;
        RECT 138.775 99.540 139.775 100.540 ;
        RECT 140.775 99.540 141.775 100.540 ;
        RECT 142.775 99.540 143.775 100.540 ;
        RECT 144.775 99.540 145.775 100.540 ;
        RECT 146.775 99.540 147.775 100.540 ;
        RECT 148.775 99.540 149.775 100.540 ;
        RECT 150.775 99.540 151.775 100.540 ;
        RECT 152.775 99.540 153.775 100.540 ;
        RECT 7.690 98.690 7.990 99.540 ;
        RECT 9.690 98.690 9.990 99.540 ;
        RECT 11.690 98.690 11.990 99.540 ;
        RECT 13.690 98.690 13.990 99.540 ;
        RECT 15.690 98.690 15.990 99.540 ;
        RECT 17.690 98.690 17.990 99.540 ;
        RECT 19.690 98.690 19.990 99.540 ;
        RECT 21.690 98.690 21.990 99.540 ;
        RECT 23.690 98.690 23.990 99.540 ;
        RECT 25.690 98.690 25.990 99.540 ;
        RECT 27.690 98.690 27.990 99.540 ;
        RECT 29.690 98.690 29.990 99.540 ;
        RECT 31.690 98.690 31.990 99.540 ;
        RECT 33.690 98.690 33.990 99.540 ;
        RECT 35.690 98.690 35.990 99.540 ;
        RECT 37.690 98.690 37.990 99.540 ;
        RECT 39.690 98.690 39.990 99.540 ;
        RECT 41.690 98.690 41.990 99.540 ;
        RECT 43.690 98.690 43.990 99.540 ;
        RECT 45.690 98.690 45.990 99.540 ;
        RECT 47.690 98.690 47.990 99.540 ;
        RECT 49.690 98.690 49.990 99.540 ;
        RECT 51.690 98.690 51.990 99.540 ;
        RECT 53.690 98.690 53.990 99.540 ;
        RECT 55.690 98.690 55.990 99.540 ;
        RECT 57.690 98.690 57.990 99.540 ;
        RECT 59.690 98.690 59.990 99.540 ;
        RECT 61.690 98.690 61.990 99.540 ;
        RECT 63.690 98.690 63.990 99.540 ;
        RECT 65.690 98.690 65.990 99.540 ;
        RECT 67.690 98.690 67.990 99.540 ;
        RECT 69.690 98.690 69.990 99.540 ;
        RECT 71.690 98.690 71.990 99.540 ;
        RECT 73.690 98.690 73.990 99.540 ;
        RECT 87.125 98.690 87.425 99.540 ;
        RECT 89.125 98.690 89.425 99.540 ;
        RECT 91.125 98.690 91.425 99.540 ;
        RECT 93.125 98.690 93.425 99.540 ;
        RECT 95.125 98.690 95.425 99.540 ;
        RECT 97.125 98.690 97.425 99.540 ;
        RECT 99.125 98.690 99.425 99.540 ;
        RECT 101.125 98.690 101.425 99.540 ;
        RECT 103.125 98.690 103.425 99.540 ;
        RECT 105.125 98.690 105.425 99.540 ;
        RECT 107.125 98.690 107.425 99.540 ;
        RECT 109.125 98.690 109.425 99.540 ;
        RECT 111.125 98.690 111.425 99.540 ;
        RECT 113.125 98.690 113.425 99.540 ;
        RECT 115.125 98.690 115.425 99.540 ;
        RECT 117.125 98.690 117.425 99.540 ;
        RECT 119.125 98.690 119.425 99.540 ;
        RECT 121.125 98.690 121.425 99.540 ;
        RECT 123.125 98.690 123.425 99.540 ;
        RECT 125.125 98.690 125.425 99.540 ;
        RECT 127.125 98.690 127.425 99.540 ;
        RECT 129.125 98.690 129.425 99.540 ;
        RECT 131.125 98.690 131.425 99.540 ;
        RECT 133.125 98.690 133.425 99.540 ;
        RECT 135.125 98.690 135.425 99.540 ;
        RECT 137.125 98.690 137.425 99.540 ;
        RECT 139.125 98.690 139.425 99.540 ;
        RECT 141.125 98.690 141.425 99.540 ;
        RECT 143.125 98.690 143.425 99.540 ;
        RECT 145.125 98.690 145.425 99.540 ;
        RECT 147.125 98.690 147.425 99.540 ;
        RECT 149.125 98.690 149.425 99.540 ;
        RECT 151.125 98.690 151.425 99.540 ;
        RECT 153.125 98.690 153.425 99.540 ;
        RECT 7.340 97.690 8.340 98.690 ;
        RECT 9.340 97.690 10.340 98.690 ;
        RECT 11.340 97.690 12.340 98.690 ;
        RECT 13.340 97.690 14.340 98.690 ;
        RECT 15.340 97.690 16.340 98.690 ;
        RECT 17.340 97.690 18.340 98.690 ;
        RECT 19.340 97.690 20.340 98.690 ;
        RECT 21.340 97.690 22.340 98.690 ;
        RECT 23.340 97.690 24.340 98.690 ;
        RECT 25.340 97.690 26.340 98.690 ;
        RECT 27.340 97.690 28.340 98.690 ;
        RECT 29.340 97.690 30.340 98.690 ;
        RECT 31.340 97.690 32.340 98.690 ;
        RECT 33.340 97.690 34.340 98.690 ;
        RECT 35.340 97.690 36.340 98.690 ;
        RECT 37.340 97.690 38.340 98.690 ;
        RECT 39.340 97.690 40.340 98.690 ;
        RECT 41.340 97.690 42.340 98.690 ;
        RECT 43.340 97.690 44.340 98.690 ;
        RECT 45.340 97.690 46.340 98.690 ;
        RECT 47.340 97.690 48.340 98.690 ;
        RECT 49.340 97.690 50.340 98.690 ;
        RECT 51.340 97.690 52.340 98.690 ;
        RECT 53.340 97.690 54.340 98.690 ;
        RECT 55.340 97.690 56.340 98.690 ;
        RECT 57.340 97.690 58.340 98.690 ;
        RECT 59.340 97.690 60.340 98.690 ;
        RECT 61.340 97.690 62.340 98.690 ;
        RECT 63.340 97.690 64.340 98.690 ;
        RECT 65.340 97.690 66.340 98.690 ;
        RECT 67.340 97.690 68.340 98.690 ;
        RECT 69.340 97.690 70.340 98.690 ;
        RECT 71.340 97.690 72.340 98.690 ;
        RECT 73.340 97.690 74.340 98.690 ;
        RECT 86.775 97.690 87.775 98.690 ;
        RECT 88.775 97.690 89.775 98.690 ;
        RECT 90.775 97.690 91.775 98.690 ;
        RECT 92.775 97.690 93.775 98.690 ;
        RECT 94.775 97.690 95.775 98.690 ;
        RECT 96.775 97.690 97.775 98.690 ;
        RECT 98.775 97.690 99.775 98.690 ;
        RECT 100.775 97.690 101.775 98.690 ;
        RECT 102.775 97.690 103.775 98.690 ;
        RECT 104.775 97.690 105.775 98.690 ;
        RECT 106.775 97.690 107.775 98.690 ;
        RECT 108.775 97.690 109.775 98.690 ;
        RECT 110.775 97.690 111.775 98.690 ;
        RECT 112.775 97.690 113.775 98.690 ;
        RECT 114.775 97.690 115.775 98.690 ;
        RECT 116.775 97.690 117.775 98.690 ;
        RECT 118.775 97.690 119.775 98.690 ;
        RECT 120.775 97.690 121.775 98.690 ;
        RECT 122.775 97.690 123.775 98.690 ;
        RECT 124.775 97.690 125.775 98.690 ;
        RECT 126.775 97.690 127.775 98.690 ;
        RECT 128.775 97.690 129.775 98.690 ;
        RECT 130.775 97.690 131.775 98.690 ;
        RECT 132.775 97.690 133.775 98.690 ;
        RECT 134.775 97.690 135.775 98.690 ;
        RECT 136.775 97.690 137.775 98.690 ;
        RECT 138.775 97.690 139.775 98.690 ;
        RECT 140.775 97.690 141.775 98.690 ;
        RECT 142.775 97.690 143.775 98.690 ;
        RECT 144.775 97.690 145.775 98.690 ;
        RECT 146.775 97.690 147.775 98.690 ;
        RECT 148.775 97.690 149.775 98.690 ;
        RECT 150.775 97.690 151.775 98.690 ;
        RECT 152.775 97.690 153.775 98.690 ;
        RECT 7.690 96.840 7.990 97.690 ;
        RECT 9.690 96.840 9.990 97.690 ;
        RECT 11.690 96.840 11.990 97.690 ;
        RECT 13.690 96.840 13.990 97.690 ;
        RECT 15.690 96.840 15.990 97.690 ;
        RECT 17.690 96.840 17.990 97.690 ;
        RECT 19.690 96.840 19.990 97.690 ;
        RECT 21.690 96.840 21.990 97.690 ;
        RECT 23.690 96.840 23.990 97.690 ;
        RECT 25.690 96.840 25.990 97.690 ;
        RECT 27.690 96.840 27.990 97.690 ;
        RECT 29.690 96.840 29.990 97.690 ;
        RECT 31.690 96.840 31.990 97.690 ;
        RECT 33.690 96.840 33.990 97.690 ;
        RECT 35.690 96.840 35.990 97.690 ;
        RECT 37.690 96.840 37.990 97.690 ;
        RECT 39.690 96.840 39.990 97.690 ;
        RECT 41.690 96.840 41.990 97.690 ;
        RECT 43.690 96.840 43.990 97.690 ;
        RECT 45.690 96.840 45.990 97.690 ;
        RECT 47.690 96.840 47.990 97.690 ;
        RECT 49.690 96.840 49.990 97.690 ;
        RECT 51.690 96.840 51.990 97.690 ;
        RECT 53.690 96.840 53.990 97.690 ;
        RECT 55.690 96.840 55.990 97.690 ;
        RECT 57.690 96.840 57.990 97.690 ;
        RECT 59.690 96.840 59.990 97.690 ;
        RECT 61.690 96.840 61.990 97.690 ;
        RECT 63.690 96.840 63.990 97.690 ;
        RECT 65.690 96.840 65.990 97.690 ;
        RECT 67.690 96.840 67.990 97.690 ;
        RECT 69.690 96.840 69.990 97.690 ;
        RECT 71.690 96.840 71.990 97.690 ;
        RECT 73.690 96.840 73.990 97.690 ;
        RECT 87.125 96.840 87.425 97.690 ;
        RECT 89.125 96.840 89.425 97.690 ;
        RECT 91.125 96.840 91.425 97.690 ;
        RECT 93.125 96.840 93.425 97.690 ;
        RECT 95.125 96.840 95.425 97.690 ;
        RECT 97.125 96.840 97.425 97.690 ;
        RECT 99.125 96.840 99.425 97.690 ;
        RECT 101.125 96.840 101.425 97.690 ;
        RECT 103.125 96.840 103.425 97.690 ;
        RECT 105.125 96.840 105.425 97.690 ;
        RECT 107.125 96.840 107.425 97.690 ;
        RECT 109.125 96.840 109.425 97.690 ;
        RECT 111.125 96.840 111.425 97.690 ;
        RECT 113.125 96.840 113.425 97.690 ;
        RECT 115.125 96.840 115.425 97.690 ;
        RECT 117.125 96.840 117.425 97.690 ;
        RECT 119.125 96.840 119.425 97.690 ;
        RECT 121.125 96.840 121.425 97.690 ;
        RECT 123.125 96.840 123.425 97.690 ;
        RECT 125.125 96.840 125.425 97.690 ;
        RECT 127.125 96.840 127.425 97.690 ;
        RECT 129.125 96.840 129.425 97.690 ;
        RECT 131.125 96.840 131.425 97.690 ;
        RECT 133.125 96.840 133.425 97.690 ;
        RECT 135.125 96.840 135.425 97.690 ;
        RECT 137.125 96.840 137.425 97.690 ;
        RECT 139.125 96.840 139.425 97.690 ;
        RECT 141.125 96.840 141.425 97.690 ;
        RECT 143.125 96.840 143.425 97.690 ;
        RECT 145.125 96.840 145.425 97.690 ;
        RECT 147.125 96.840 147.425 97.690 ;
        RECT 149.125 96.840 149.425 97.690 ;
        RECT 151.125 96.840 151.425 97.690 ;
        RECT 153.125 96.840 153.425 97.690 ;
        RECT 7.340 95.840 8.340 96.840 ;
        RECT 9.340 95.840 10.340 96.840 ;
        RECT 11.340 95.840 12.340 96.840 ;
        RECT 13.340 95.840 14.340 96.840 ;
        RECT 15.340 95.840 16.340 96.840 ;
        RECT 17.340 95.840 18.340 96.840 ;
        RECT 19.340 95.840 20.340 96.840 ;
        RECT 21.340 95.840 22.340 96.840 ;
        RECT 23.340 95.840 24.340 96.840 ;
        RECT 25.340 95.840 26.340 96.840 ;
        RECT 27.340 95.840 28.340 96.840 ;
        RECT 29.340 95.840 30.340 96.840 ;
        RECT 31.340 95.840 32.340 96.840 ;
        RECT 33.340 95.840 34.340 96.840 ;
        RECT 35.340 95.840 36.340 96.840 ;
        RECT 37.340 95.840 38.340 96.840 ;
        RECT 39.340 95.840 40.340 96.840 ;
        RECT 41.340 95.840 42.340 96.840 ;
        RECT 43.340 95.840 44.340 96.840 ;
        RECT 45.340 95.840 46.340 96.840 ;
        RECT 47.340 95.840 48.340 96.840 ;
        RECT 49.340 95.840 50.340 96.840 ;
        RECT 51.340 95.840 52.340 96.840 ;
        RECT 53.340 95.840 54.340 96.840 ;
        RECT 55.340 95.840 56.340 96.840 ;
        RECT 57.340 95.840 58.340 96.840 ;
        RECT 59.340 95.840 60.340 96.840 ;
        RECT 61.340 95.840 62.340 96.840 ;
        RECT 63.340 95.840 64.340 96.840 ;
        RECT 65.340 95.840 66.340 96.840 ;
        RECT 67.340 95.840 68.340 96.840 ;
        RECT 69.340 95.840 70.340 96.840 ;
        RECT 71.340 95.840 72.340 96.840 ;
        RECT 73.340 95.840 74.340 96.840 ;
        RECT 86.775 95.840 87.775 96.840 ;
        RECT 88.775 95.840 89.775 96.840 ;
        RECT 90.775 95.840 91.775 96.840 ;
        RECT 92.775 95.840 93.775 96.840 ;
        RECT 94.775 95.840 95.775 96.840 ;
        RECT 96.775 95.840 97.775 96.840 ;
        RECT 98.775 95.840 99.775 96.840 ;
        RECT 100.775 95.840 101.775 96.840 ;
        RECT 102.775 95.840 103.775 96.840 ;
        RECT 104.775 95.840 105.775 96.840 ;
        RECT 106.775 95.840 107.775 96.840 ;
        RECT 108.775 95.840 109.775 96.840 ;
        RECT 110.775 95.840 111.775 96.840 ;
        RECT 112.775 95.840 113.775 96.840 ;
        RECT 114.775 95.840 115.775 96.840 ;
        RECT 116.775 95.840 117.775 96.840 ;
        RECT 118.775 95.840 119.775 96.840 ;
        RECT 120.775 95.840 121.775 96.840 ;
        RECT 122.775 95.840 123.775 96.840 ;
        RECT 124.775 95.840 125.775 96.840 ;
        RECT 126.775 95.840 127.775 96.840 ;
        RECT 128.775 95.840 129.775 96.840 ;
        RECT 130.775 95.840 131.775 96.840 ;
        RECT 132.775 95.840 133.775 96.840 ;
        RECT 134.775 95.840 135.775 96.840 ;
        RECT 136.775 95.840 137.775 96.840 ;
        RECT 138.775 95.840 139.775 96.840 ;
        RECT 140.775 95.840 141.775 96.840 ;
        RECT 142.775 95.840 143.775 96.840 ;
        RECT 144.775 95.840 145.775 96.840 ;
        RECT 146.775 95.840 147.775 96.840 ;
        RECT 148.775 95.840 149.775 96.840 ;
        RECT 150.775 95.840 151.775 96.840 ;
        RECT 152.775 95.840 153.775 96.840 ;
        RECT 7.690 94.990 7.990 95.840 ;
        RECT 9.690 94.990 9.990 95.840 ;
        RECT 11.690 94.990 11.990 95.840 ;
        RECT 13.690 94.990 13.990 95.840 ;
        RECT 15.690 94.990 15.990 95.840 ;
        RECT 17.690 94.990 17.990 95.840 ;
        RECT 19.690 94.990 19.990 95.840 ;
        RECT 21.690 94.990 21.990 95.840 ;
        RECT 23.690 94.990 23.990 95.840 ;
        RECT 25.690 94.990 25.990 95.840 ;
        RECT 27.690 94.990 27.990 95.840 ;
        RECT 29.690 94.990 29.990 95.840 ;
        RECT 31.690 94.990 31.990 95.840 ;
        RECT 33.690 94.990 33.990 95.840 ;
        RECT 35.690 94.990 35.990 95.840 ;
        RECT 37.690 94.990 37.990 95.840 ;
        RECT 39.690 94.990 39.990 95.840 ;
        RECT 41.690 94.990 41.990 95.840 ;
        RECT 43.690 94.990 43.990 95.840 ;
        RECT 45.690 94.990 45.990 95.840 ;
        RECT 47.690 94.990 47.990 95.840 ;
        RECT 49.690 94.990 49.990 95.840 ;
        RECT 51.690 94.990 51.990 95.840 ;
        RECT 53.690 94.990 53.990 95.840 ;
        RECT 55.690 94.990 55.990 95.840 ;
        RECT 57.690 94.990 57.990 95.840 ;
        RECT 59.690 94.990 59.990 95.840 ;
        RECT 61.690 94.990 61.990 95.840 ;
        RECT 63.690 94.990 63.990 95.840 ;
        RECT 65.690 94.990 65.990 95.840 ;
        RECT 67.690 94.990 67.990 95.840 ;
        RECT 69.690 94.990 69.990 95.840 ;
        RECT 71.690 94.990 71.990 95.840 ;
        RECT 73.690 94.990 73.990 95.840 ;
        RECT 87.125 94.990 87.425 95.840 ;
        RECT 89.125 94.990 89.425 95.840 ;
        RECT 91.125 94.990 91.425 95.840 ;
        RECT 93.125 94.990 93.425 95.840 ;
        RECT 95.125 94.990 95.425 95.840 ;
        RECT 97.125 94.990 97.425 95.840 ;
        RECT 99.125 94.990 99.425 95.840 ;
        RECT 101.125 94.990 101.425 95.840 ;
        RECT 103.125 94.990 103.425 95.840 ;
        RECT 105.125 94.990 105.425 95.840 ;
        RECT 107.125 94.990 107.425 95.840 ;
        RECT 109.125 94.990 109.425 95.840 ;
        RECT 111.125 94.990 111.425 95.840 ;
        RECT 113.125 94.990 113.425 95.840 ;
        RECT 115.125 94.990 115.425 95.840 ;
        RECT 117.125 94.990 117.425 95.840 ;
        RECT 119.125 94.990 119.425 95.840 ;
        RECT 121.125 94.990 121.425 95.840 ;
        RECT 123.125 94.990 123.425 95.840 ;
        RECT 125.125 94.990 125.425 95.840 ;
        RECT 127.125 94.990 127.425 95.840 ;
        RECT 129.125 94.990 129.425 95.840 ;
        RECT 131.125 94.990 131.425 95.840 ;
        RECT 133.125 94.990 133.425 95.840 ;
        RECT 135.125 94.990 135.425 95.840 ;
        RECT 137.125 94.990 137.425 95.840 ;
        RECT 139.125 94.990 139.425 95.840 ;
        RECT 141.125 94.990 141.425 95.840 ;
        RECT 143.125 94.990 143.425 95.840 ;
        RECT 145.125 94.990 145.425 95.840 ;
        RECT 147.125 94.990 147.425 95.840 ;
        RECT 149.125 94.990 149.425 95.840 ;
        RECT 151.125 94.990 151.425 95.840 ;
        RECT 153.125 94.990 153.425 95.840 ;
        RECT 7.340 93.990 8.340 94.990 ;
        RECT 9.340 93.990 10.340 94.990 ;
        RECT 11.340 93.990 12.340 94.990 ;
        RECT 13.340 93.990 14.340 94.990 ;
        RECT 15.340 93.990 16.340 94.990 ;
        RECT 17.340 93.990 18.340 94.990 ;
        RECT 19.340 93.990 20.340 94.990 ;
        RECT 21.340 93.990 22.340 94.990 ;
        RECT 23.340 93.990 24.340 94.990 ;
        RECT 25.340 93.990 26.340 94.990 ;
        RECT 27.340 93.990 28.340 94.990 ;
        RECT 29.340 93.990 30.340 94.990 ;
        RECT 31.340 93.990 32.340 94.990 ;
        RECT 33.340 93.990 34.340 94.990 ;
        RECT 35.340 93.990 36.340 94.990 ;
        RECT 37.340 93.990 38.340 94.990 ;
        RECT 39.340 93.990 40.340 94.990 ;
        RECT 41.340 93.990 42.340 94.990 ;
        RECT 43.340 93.990 44.340 94.990 ;
        RECT 45.340 93.990 46.340 94.990 ;
        RECT 47.340 93.990 48.340 94.990 ;
        RECT 49.340 93.990 50.340 94.990 ;
        RECT 51.340 93.990 52.340 94.990 ;
        RECT 53.340 93.990 54.340 94.990 ;
        RECT 55.340 93.990 56.340 94.990 ;
        RECT 57.340 93.990 58.340 94.990 ;
        RECT 59.340 93.990 60.340 94.990 ;
        RECT 61.340 93.990 62.340 94.990 ;
        RECT 63.340 93.990 64.340 94.990 ;
        RECT 65.340 93.990 66.340 94.990 ;
        RECT 67.340 93.990 68.340 94.990 ;
        RECT 69.340 93.990 70.340 94.990 ;
        RECT 71.340 93.990 72.340 94.990 ;
        RECT 73.340 93.990 74.340 94.990 ;
        RECT 86.775 93.990 87.775 94.990 ;
        RECT 88.775 93.990 89.775 94.990 ;
        RECT 90.775 93.990 91.775 94.990 ;
        RECT 92.775 93.990 93.775 94.990 ;
        RECT 94.775 93.990 95.775 94.990 ;
        RECT 96.775 93.990 97.775 94.990 ;
        RECT 98.775 93.990 99.775 94.990 ;
        RECT 100.775 93.990 101.775 94.990 ;
        RECT 102.775 93.990 103.775 94.990 ;
        RECT 104.775 93.990 105.775 94.990 ;
        RECT 106.775 93.990 107.775 94.990 ;
        RECT 108.775 93.990 109.775 94.990 ;
        RECT 110.775 93.990 111.775 94.990 ;
        RECT 112.775 93.990 113.775 94.990 ;
        RECT 114.775 93.990 115.775 94.990 ;
        RECT 116.775 93.990 117.775 94.990 ;
        RECT 118.775 93.990 119.775 94.990 ;
        RECT 120.775 93.990 121.775 94.990 ;
        RECT 122.775 93.990 123.775 94.990 ;
        RECT 124.775 93.990 125.775 94.990 ;
        RECT 126.775 93.990 127.775 94.990 ;
        RECT 128.775 93.990 129.775 94.990 ;
        RECT 130.775 93.990 131.775 94.990 ;
        RECT 132.775 93.990 133.775 94.990 ;
        RECT 134.775 93.990 135.775 94.990 ;
        RECT 136.775 93.990 137.775 94.990 ;
        RECT 138.775 93.990 139.775 94.990 ;
        RECT 140.775 93.990 141.775 94.990 ;
        RECT 142.775 93.990 143.775 94.990 ;
        RECT 144.775 93.990 145.775 94.990 ;
        RECT 146.775 93.990 147.775 94.990 ;
        RECT 148.775 93.990 149.775 94.990 ;
        RECT 150.775 93.990 151.775 94.990 ;
        RECT 152.775 93.990 153.775 94.990 ;
        RECT 7.690 93.140 7.990 93.990 ;
        RECT 9.690 93.140 9.990 93.990 ;
        RECT 11.690 93.140 11.990 93.990 ;
        RECT 13.690 93.140 13.990 93.990 ;
        RECT 15.690 93.140 15.990 93.990 ;
        RECT 17.690 93.140 17.990 93.990 ;
        RECT 19.690 93.140 19.990 93.990 ;
        RECT 21.690 93.140 21.990 93.990 ;
        RECT 23.690 93.140 23.990 93.990 ;
        RECT 25.690 93.140 25.990 93.990 ;
        RECT 27.690 93.140 27.990 93.990 ;
        RECT 29.690 93.140 29.990 93.990 ;
        RECT 31.690 93.140 31.990 93.990 ;
        RECT 33.690 93.140 33.990 93.990 ;
        RECT 35.690 93.140 35.990 93.990 ;
        RECT 37.690 93.140 37.990 93.990 ;
        RECT 39.690 93.140 39.990 93.990 ;
        RECT 41.690 93.140 41.990 93.990 ;
        RECT 43.690 93.140 43.990 93.990 ;
        RECT 45.690 93.140 45.990 93.990 ;
        RECT 47.690 93.140 47.990 93.990 ;
        RECT 49.690 93.140 49.990 93.990 ;
        RECT 51.690 93.140 51.990 93.990 ;
        RECT 53.690 93.140 53.990 93.990 ;
        RECT 55.690 93.140 55.990 93.990 ;
        RECT 57.690 93.140 57.990 93.990 ;
        RECT 59.690 93.140 59.990 93.990 ;
        RECT 61.690 93.140 61.990 93.990 ;
        RECT 63.690 93.140 63.990 93.990 ;
        RECT 65.690 93.140 65.990 93.990 ;
        RECT 67.690 93.140 67.990 93.990 ;
        RECT 69.690 93.140 69.990 93.990 ;
        RECT 71.690 93.140 71.990 93.990 ;
        RECT 73.690 93.140 73.990 93.990 ;
        RECT 87.125 93.140 87.425 93.990 ;
        RECT 89.125 93.140 89.425 93.990 ;
        RECT 91.125 93.140 91.425 93.990 ;
        RECT 93.125 93.140 93.425 93.990 ;
        RECT 95.125 93.140 95.425 93.990 ;
        RECT 97.125 93.140 97.425 93.990 ;
        RECT 99.125 93.140 99.425 93.990 ;
        RECT 101.125 93.140 101.425 93.990 ;
        RECT 103.125 93.140 103.425 93.990 ;
        RECT 105.125 93.140 105.425 93.990 ;
        RECT 107.125 93.140 107.425 93.990 ;
        RECT 109.125 93.140 109.425 93.990 ;
        RECT 111.125 93.140 111.425 93.990 ;
        RECT 113.125 93.140 113.425 93.990 ;
        RECT 115.125 93.140 115.425 93.990 ;
        RECT 117.125 93.140 117.425 93.990 ;
        RECT 119.125 93.140 119.425 93.990 ;
        RECT 121.125 93.140 121.425 93.990 ;
        RECT 123.125 93.140 123.425 93.990 ;
        RECT 125.125 93.140 125.425 93.990 ;
        RECT 127.125 93.140 127.425 93.990 ;
        RECT 129.125 93.140 129.425 93.990 ;
        RECT 131.125 93.140 131.425 93.990 ;
        RECT 133.125 93.140 133.425 93.990 ;
        RECT 135.125 93.140 135.425 93.990 ;
        RECT 137.125 93.140 137.425 93.990 ;
        RECT 139.125 93.140 139.425 93.990 ;
        RECT 141.125 93.140 141.425 93.990 ;
        RECT 143.125 93.140 143.425 93.990 ;
        RECT 145.125 93.140 145.425 93.990 ;
        RECT 147.125 93.140 147.425 93.990 ;
        RECT 149.125 93.140 149.425 93.990 ;
        RECT 151.125 93.140 151.425 93.990 ;
        RECT 153.125 93.140 153.425 93.990 ;
        RECT 7.340 92.140 8.340 93.140 ;
        RECT 9.340 92.140 10.340 93.140 ;
        RECT 11.340 92.140 12.340 93.140 ;
        RECT 13.340 92.140 14.340 93.140 ;
        RECT 15.340 92.140 16.340 93.140 ;
        RECT 17.340 92.140 18.340 93.140 ;
        RECT 19.340 92.140 20.340 93.140 ;
        RECT 21.340 92.140 22.340 93.140 ;
        RECT 23.340 92.140 24.340 93.140 ;
        RECT 25.340 92.140 26.340 93.140 ;
        RECT 27.340 92.140 28.340 93.140 ;
        RECT 29.340 92.140 30.340 93.140 ;
        RECT 31.340 92.140 32.340 93.140 ;
        RECT 33.340 92.140 34.340 93.140 ;
        RECT 35.340 92.140 36.340 93.140 ;
        RECT 37.340 92.140 38.340 93.140 ;
        RECT 39.340 92.140 40.340 93.140 ;
        RECT 41.340 92.140 42.340 93.140 ;
        RECT 43.340 92.140 44.340 93.140 ;
        RECT 45.340 92.140 46.340 93.140 ;
        RECT 47.340 92.140 48.340 93.140 ;
        RECT 49.340 92.140 50.340 93.140 ;
        RECT 51.340 92.140 52.340 93.140 ;
        RECT 53.340 92.140 54.340 93.140 ;
        RECT 55.340 92.140 56.340 93.140 ;
        RECT 57.340 92.140 58.340 93.140 ;
        RECT 59.340 92.140 60.340 93.140 ;
        RECT 61.340 92.140 62.340 93.140 ;
        RECT 63.340 92.140 64.340 93.140 ;
        RECT 65.340 92.140 66.340 93.140 ;
        RECT 67.340 92.140 68.340 93.140 ;
        RECT 69.340 92.140 70.340 93.140 ;
        RECT 71.340 92.140 72.340 93.140 ;
        RECT 73.340 92.140 74.340 93.140 ;
        RECT 86.775 92.140 87.775 93.140 ;
        RECT 88.775 92.140 89.775 93.140 ;
        RECT 90.775 92.140 91.775 93.140 ;
        RECT 92.775 92.140 93.775 93.140 ;
        RECT 94.775 92.140 95.775 93.140 ;
        RECT 96.775 92.140 97.775 93.140 ;
        RECT 98.775 92.140 99.775 93.140 ;
        RECT 100.775 92.140 101.775 93.140 ;
        RECT 102.775 92.140 103.775 93.140 ;
        RECT 104.775 92.140 105.775 93.140 ;
        RECT 106.775 92.140 107.775 93.140 ;
        RECT 108.775 92.140 109.775 93.140 ;
        RECT 110.775 92.140 111.775 93.140 ;
        RECT 112.775 92.140 113.775 93.140 ;
        RECT 114.775 92.140 115.775 93.140 ;
        RECT 116.775 92.140 117.775 93.140 ;
        RECT 118.775 92.140 119.775 93.140 ;
        RECT 120.775 92.140 121.775 93.140 ;
        RECT 122.775 92.140 123.775 93.140 ;
        RECT 124.775 92.140 125.775 93.140 ;
        RECT 126.775 92.140 127.775 93.140 ;
        RECT 128.775 92.140 129.775 93.140 ;
        RECT 130.775 92.140 131.775 93.140 ;
        RECT 132.775 92.140 133.775 93.140 ;
        RECT 134.775 92.140 135.775 93.140 ;
        RECT 136.775 92.140 137.775 93.140 ;
        RECT 138.775 92.140 139.775 93.140 ;
        RECT 140.775 92.140 141.775 93.140 ;
        RECT 142.775 92.140 143.775 93.140 ;
        RECT 144.775 92.140 145.775 93.140 ;
        RECT 146.775 92.140 147.775 93.140 ;
        RECT 148.775 92.140 149.775 93.140 ;
        RECT 150.775 92.140 151.775 93.140 ;
        RECT 152.775 92.140 153.775 93.140 ;
        RECT 7.690 91.290 7.990 92.140 ;
        RECT 9.690 91.290 9.990 92.140 ;
        RECT 11.690 91.290 11.990 92.140 ;
        RECT 13.690 91.290 13.990 92.140 ;
        RECT 15.690 91.290 15.990 92.140 ;
        RECT 17.690 91.290 17.990 92.140 ;
        RECT 19.690 91.290 19.990 92.140 ;
        RECT 21.690 91.290 21.990 92.140 ;
        RECT 23.690 91.290 23.990 92.140 ;
        RECT 25.690 91.290 25.990 92.140 ;
        RECT 27.690 91.290 27.990 92.140 ;
        RECT 29.690 91.290 29.990 92.140 ;
        RECT 31.690 91.290 31.990 92.140 ;
        RECT 33.690 91.290 33.990 92.140 ;
        RECT 35.690 91.290 35.990 92.140 ;
        RECT 37.690 91.290 37.990 92.140 ;
        RECT 39.690 91.290 39.990 92.140 ;
        RECT 41.690 91.290 41.990 92.140 ;
        RECT 43.690 91.290 43.990 92.140 ;
        RECT 45.690 91.290 45.990 92.140 ;
        RECT 47.690 91.290 47.990 92.140 ;
        RECT 49.690 91.290 49.990 92.140 ;
        RECT 51.690 91.290 51.990 92.140 ;
        RECT 53.690 91.290 53.990 92.140 ;
        RECT 55.690 91.290 55.990 92.140 ;
        RECT 57.690 91.290 57.990 92.140 ;
        RECT 59.690 91.290 59.990 92.140 ;
        RECT 61.690 91.290 61.990 92.140 ;
        RECT 63.690 91.290 63.990 92.140 ;
        RECT 65.690 91.290 65.990 92.140 ;
        RECT 67.690 91.290 67.990 92.140 ;
        RECT 69.690 91.290 69.990 92.140 ;
        RECT 71.690 91.290 71.990 92.140 ;
        RECT 73.690 91.290 73.990 92.140 ;
        RECT 87.125 91.290 87.425 92.140 ;
        RECT 89.125 91.290 89.425 92.140 ;
        RECT 91.125 91.290 91.425 92.140 ;
        RECT 93.125 91.290 93.425 92.140 ;
        RECT 95.125 91.290 95.425 92.140 ;
        RECT 97.125 91.290 97.425 92.140 ;
        RECT 99.125 91.290 99.425 92.140 ;
        RECT 101.125 91.290 101.425 92.140 ;
        RECT 103.125 91.290 103.425 92.140 ;
        RECT 105.125 91.290 105.425 92.140 ;
        RECT 107.125 91.290 107.425 92.140 ;
        RECT 109.125 91.290 109.425 92.140 ;
        RECT 111.125 91.290 111.425 92.140 ;
        RECT 113.125 91.290 113.425 92.140 ;
        RECT 115.125 91.290 115.425 92.140 ;
        RECT 117.125 91.290 117.425 92.140 ;
        RECT 119.125 91.290 119.425 92.140 ;
        RECT 121.125 91.290 121.425 92.140 ;
        RECT 123.125 91.290 123.425 92.140 ;
        RECT 125.125 91.290 125.425 92.140 ;
        RECT 127.125 91.290 127.425 92.140 ;
        RECT 129.125 91.290 129.425 92.140 ;
        RECT 131.125 91.290 131.425 92.140 ;
        RECT 133.125 91.290 133.425 92.140 ;
        RECT 135.125 91.290 135.425 92.140 ;
        RECT 137.125 91.290 137.425 92.140 ;
        RECT 139.125 91.290 139.425 92.140 ;
        RECT 141.125 91.290 141.425 92.140 ;
        RECT 143.125 91.290 143.425 92.140 ;
        RECT 145.125 91.290 145.425 92.140 ;
        RECT 147.125 91.290 147.425 92.140 ;
        RECT 149.125 91.290 149.425 92.140 ;
        RECT 151.125 91.290 151.425 92.140 ;
        RECT 153.125 91.290 153.425 92.140 ;
        RECT 7.340 90.290 8.340 91.290 ;
        RECT 9.340 90.290 10.340 91.290 ;
        RECT 11.340 90.290 12.340 91.290 ;
        RECT 13.340 90.290 14.340 91.290 ;
        RECT 15.340 90.290 16.340 91.290 ;
        RECT 17.340 90.290 18.340 91.290 ;
        RECT 19.340 90.290 20.340 91.290 ;
        RECT 21.340 90.290 22.340 91.290 ;
        RECT 23.340 90.290 24.340 91.290 ;
        RECT 25.340 90.290 26.340 91.290 ;
        RECT 27.340 90.290 28.340 91.290 ;
        RECT 29.340 90.290 30.340 91.290 ;
        RECT 31.340 90.290 32.340 91.290 ;
        RECT 33.340 90.290 34.340 91.290 ;
        RECT 35.340 90.290 36.340 91.290 ;
        RECT 37.340 90.290 38.340 91.290 ;
        RECT 39.340 90.290 40.340 91.290 ;
        RECT 41.340 90.290 42.340 91.290 ;
        RECT 43.340 90.290 44.340 91.290 ;
        RECT 45.340 90.290 46.340 91.290 ;
        RECT 47.340 90.290 48.340 91.290 ;
        RECT 49.340 90.290 50.340 91.290 ;
        RECT 51.340 90.290 52.340 91.290 ;
        RECT 53.340 90.290 54.340 91.290 ;
        RECT 55.340 90.290 56.340 91.290 ;
        RECT 57.340 90.290 58.340 91.290 ;
        RECT 59.340 90.290 60.340 91.290 ;
        RECT 61.340 90.290 62.340 91.290 ;
        RECT 63.340 90.290 64.340 91.290 ;
        RECT 65.340 90.290 66.340 91.290 ;
        RECT 67.340 90.290 68.340 91.290 ;
        RECT 69.340 90.290 70.340 91.290 ;
        RECT 71.340 90.290 72.340 91.290 ;
        RECT 73.340 90.290 74.340 91.290 ;
        RECT 86.775 90.290 87.775 91.290 ;
        RECT 88.775 90.290 89.775 91.290 ;
        RECT 90.775 90.290 91.775 91.290 ;
        RECT 92.775 90.290 93.775 91.290 ;
        RECT 94.775 90.290 95.775 91.290 ;
        RECT 96.775 90.290 97.775 91.290 ;
        RECT 98.775 90.290 99.775 91.290 ;
        RECT 100.775 90.290 101.775 91.290 ;
        RECT 102.775 90.290 103.775 91.290 ;
        RECT 104.775 90.290 105.775 91.290 ;
        RECT 106.775 90.290 107.775 91.290 ;
        RECT 108.775 90.290 109.775 91.290 ;
        RECT 110.775 90.290 111.775 91.290 ;
        RECT 112.775 90.290 113.775 91.290 ;
        RECT 114.775 90.290 115.775 91.290 ;
        RECT 116.775 90.290 117.775 91.290 ;
        RECT 118.775 90.290 119.775 91.290 ;
        RECT 120.775 90.290 121.775 91.290 ;
        RECT 122.775 90.290 123.775 91.290 ;
        RECT 124.775 90.290 125.775 91.290 ;
        RECT 126.775 90.290 127.775 91.290 ;
        RECT 128.775 90.290 129.775 91.290 ;
        RECT 130.775 90.290 131.775 91.290 ;
        RECT 132.775 90.290 133.775 91.290 ;
        RECT 134.775 90.290 135.775 91.290 ;
        RECT 136.775 90.290 137.775 91.290 ;
        RECT 138.775 90.290 139.775 91.290 ;
        RECT 140.775 90.290 141.775 91.290 ;
        RECT 142.775 90.290 143.775 91.290 ;
        RECT 144.775 90.290 145.775 91.290 ;
        RECT 146.775 90.290 147.775 91.290 ;
        RECT 148.775 90.290 149.775 91.290 ;
        RECT 150.775 90.290 151.775 91.290 ;
        RECT 152.775 90.290 153.775 91.290 ;
        RECT 7.690 89.440 7.990 90.290 ;
        RECT 9.690 89.440 9.990 90.290 ;
        RECT 11.690 89.440 11.990 90.290 ;
        RECT 13.690 89.440 13.990 90.290 ;
        RECT 15.690 89.440 15.990 90.290 ;
        RECT 17.690 89.440 17.990 90.290 ;
        RECT 19.690 89.440 19.990 90.290 ;
        RECT 21.690 89.440 21.990 90.290 ;
        RECT 23.690 89.440 23.990 90.290 ;
        RECT 25.690 89.440 25.990 90.290 ;
        RECT 27.690 89.440 27.990 90.290 ;
        RECT 29.690 89.440 29.990 90.290 ;
        RECT 31.690 89.440 31.990 90.290 ;
        RECT 33.690 89.440 33.990 90.290 ;
        RECT 35.690 89.440 35.990 90.290 ;
        RECT 37.690 89.440 37.990 90.290 ;
        RECT 39.690 89.440 39.990 90.290 ;
        RECT 41.690 89.440 41.990 90.290 ;
        RECT 43.690 89.440 43.990 90.290 ;
        RECT 45.690 89.440 45.990 90.290 ;
        RECT 47.690 89.440 47.990 90.290 ;
        RECT 49.690 89.440 49.990 90.290 ;
        RECT 51.690 89.440 51.990 90.290 ;
        RECT 53.690 89.440 53.990 90.290 ;
        RECT 55.690 89.440 55.990 90.290 ;
        RECT 57.690 89.440 57.990 90.290 ;
        RECT 59.690 89.440 59.990 90.290 ;
        RECT 61.690 89.440 61.990 90.290 ;
        RECT 63.690 89.440 63.990 90.290 ;
        RECT 65.690 89.440 65.990 90.290 ;
        RECT 67.690 89.440 67.990 90.290 ;
        RECT 69.690 89.440 69.990 90.290 ;
        RECT 71.690 89.440 71.990 90.290 ;
        RECT 73.690 89.440 73.990 90.290 ;
        RECT 87.125 89.440 87.425 90.290 ;
        RECT 89.125 89.440 89.425 90.290 ;
        RECT 91.125 89.440 91.425 90.290 ;
        RECT 93.125 89.440 93.425 90.290 ;
        RECT 95.125 89.440 95.425 90.290 ;
        RECT 97.125 89.440 97.425 90.290 ;
        RECT 99.125 89.440 99.425 90.290 ;
        RECT 101.125 89.440 101.425 90.290 ;
        RECT 103.125 89.440 103.425 90.290 ;
        RECT 105.125 89.440 105.425 90.290 ;
        RECT 107.125 89.440 107.425 90.290 ;
        RECT 109.125 89.440 109.425 90.290 ;
        RECT 111.125 89.440 111.425 90.290 ;
        RECT 113.125 89.440 113.425 90.290 ;
        RECT 115.125 89.440 115.425 90.290 ;
        RECT 117.125 89.440 117.425 90.290 ;
        RECT 119.125 89.440 119.425 90.290 ;
        RECT 121.125 89.440 121.425 90.290 ;
        RECT 123.125 89.440 123.425 90.290 ;
        RECT 125.125 89.440 125.425 90.290 ;
        RECT 127.125 89.440 127.425 90.290 ;
        RECT 129.125 89.440 129.425 90.290 ;
        RECT 131.125 89.440 131.425 90.290 ;
        RECT 133.125 89.440 133.425 90.290 ;
        RECT 135.125 89.440 135.425 90.290 ;
        RECT 137.125 89.440 137.425 90.290 ;
        RECT 139.125 89.440 139.425 90.290 ;
        RECT 141.125 89.440 141.425 90.290 ;
        RECT 143.125 89.440 143.425 90.290 ;
        RECT 145.125 89.440 145.425 90.290 ;
        RECT 147.125 89.440 147.425 90.290 ;
        RECT 149.125 89.440 149.425 90.290 ;
        RECT 151.125 89.440 151.425 90.290 ;
        RECT 153.125 89.440 153.425 90.290 ;
        RECT 7.340 88.440 8.340 89.440 ;
        RECT 9.340 88.440 10.340 89.440 ;
        RECT 11.340 88.440 12.340 89.440 ;
        RECT 13.340 88.440 14.340 89.440 ;
        RECT 15.340 88.440 16.340 89.440 ;
        RECT 17.340 88.440 18.340 89.440 ;
        RECT 19.340 88.440 20.340 89.440 ;
        RECT 21.340 88.440 22.340 89.440 ;
        RECT 23.340 88.440 24.340 89.440 ;
        RECT 25.340 88.440 26.340 89.440 ;
        RECT 27.340 88.440 28.340 89.440 ;
        RECT 29.340 88.440 30.340 89.440 ;
        RECT 31.340 88.440 32.340 89.440 ;
        RECT 33.340 88.440 34.340 89.440 ;
        RECT 35.340 88.440 36.340 89.440 ;
        RECT 37.340 88.440 38.340 89.440 ;
        RECT 39.340 88.440 40.340 89.440 ;
        RECT 41.340 88.440 42.340 89.440 ;
        RECT 43.340 88.440 44.340 89.440 ;
        RECT 45.340 88.440 46.340 89.440 ;
        RECT 47.340 88.440 48.340 89.440 ;
        RECT 49.340 88.440 50.340 89.440 ;
        RECT 51.340 88.440 52.340 89.440 ;
        RECT 53.340 88.440 54.340 89.440 ;
        RECT 55.340 88.440 56.340 89.440 ;
        RECT 57.340 88.440 58.340 89.440 ;
        RECT 59.340 88.440 60.340 89.440 ;
        RECT 61.340 88.440 62.340 89.440 ;
        RECT 63.340 88.440 64.340 89.440 ;
        RECT 65.340 88.440 66.340 89.440 ;
        RECT 67.340 88.440 68.340 89.440 ;
        RECT 69.340 88.440 70.340 89.440 ;
        RECT 71.340 88.440 72.340 89.440 ;
        RECT 73.340 88.440 74.340 89.440 ;
        RECT 86.775 88.440 87.775 89.440 ;
        RECT 88.775 88.440 89.775 89.440 ;
        RECT 90.775 88.440 91.775 89.440 ;
        RECT 92.775 88.440 93.775 89.440 ;
        RECT 94.775 88.440 95.775 89.440 ;
        RECT 96.775 88.440 97.775 89.440 ;
        RECT 98.775 88.440 99.775 89.440 ;
        RECT 100.775 88.440 101.775 89.440 ;
        RECT 102.775 88.440 103.775 89.440 ;
        RECT 104.775 88.440 105.775 89.440 ;
        RECT 106.775 88.440 107.775 89.440 ;
        RECT 108.775 88.440 109.775 89.440 ;
        RECT 110.775 88.440 111.775 89.440 ;
        RECT 112.775 88.440 113.775 89.440 ;
        RECT 114.775 88.440 115.775 89.440 ;
        RECT 116.775 88.440 117.775 89.440 ;
        RECT 118.775 88.440 119.775 89.440 ;
        RECT 120.775 88.440 121.775 89.440 ;
        RECT 122.775 88.440 123.775 89.440 ;
        RECT 124.775 88.440 125.775 89.440 ;
        RECT 126.775 88.440 127.775 89.440 ;
        RECT 128.775 88.440 129.775 89.440 ;
        RECT 130.775 88.440 131.775 89.440 ;
        RECT 132.775 88.440 133.775 89.440 ;
        RECT 134.775 88.440 135.775 89.440 ;
        RECT 136.775 88.440 137.775 89.440 ;
        RECT 138.775 88.440 139.775 89.440 ;
        RECT 140.775 88.440 141.775 89.440 ;
        RECT 142.775 88.440 143.775 89.440 ;
        RECT 144.775 88.440 145.775 89.440 ;
        RECT 146.775 88.440 147.775 89.440 ;
        RECT 148.775 88.440 149.775 89.440 ;
        RECT 150.775 88.440 151.775 89.440 ;
        RECT 152.775 88.440 153.775 89.440 ;
        RECT 7.690 87.590 7.990 88.440 ;
        RECT 9.690 87.590 9.990 88.440 ;
        RECT 11.690 87.590 11.990 88.440 ;
        RECT 13.690 87.590 13.990 88.440 ;
        RECT 15.690 87.590 15.990 88.440 ;
        RECT 17.690 87.590 17.990 88.440 ;
        RECT 19.690 87.590 19.990 88.440 ;
        RECT 21.690 87.590 21.990 88.440 ;
        RECT 23.690 87.590 23.990 88.440 ;
        RECT 25.690 87.590 25.990 88.440 ;
        RECT 27.690 87.590 27.990 88.440 ;
        RECT 29.690 87.590 29.990 88.440 ;
        RECT 31.690 87.590 31.990 88.440 ;
        RECT 33.690 87.590 33.990 88.440 ;
        RECT 35.690 87.590 35.990 88.440 ;
        RECT 37.690 87.590 37.990 88.440 ;
        RECT 39.690 87.590 39.990 88.440 ;
        RECT 41.690 87.590 41.990 88.440 ;
        RECT 43.690 87.590 43.990 88.440 ;
        RECT 45.690 87.590 45.990 88.440 ;
        RECT 47.690 87.590 47.990 88.440 ;
        RECT 49.690 87.590 49.990 88.440 ;
        RECT 51.690 87.590 51.990 88.440 ;
        RECT 53.690 87.590 53.990 88.440 ;
        RECT 55.690 87.590 55.990 88.440 ;
        RECT 57.690 87.590 57.990 88.440 ;
        RECT 59.690 87.590 59.990 88.440 ;
        RECT 61.690 87.590 61.990 88.440 ;
        RECT 63.690 87.590 63.990 88.440 ;
        RECT 65.690 87.590 65.990 88.440 ;
        RECT 67.690 87.590 67.990 88.440 ;
        RECT 69.690 87.590 69.990 88.440 ;
        RECT 71.690 87.590 71.990 88.440 ;
        RECT 73.690 87.590 73.990 88.440 ;
        RECT 87.125 87.590 87.425 88.440 ;
        RECT 89.125 87.590 89.425 88.440 ;
        RECT 91.125 87.590 91.425 88.440 ;
        RECT 93.125 87.590 93.425 88.440 ;
        RECT 95.125 87.590 95.425 88.440 ;
        RECT 97.125 87.590 97.425 88.440 ;
        RECT 99.125 87.590 99.425 88.440 ;
        RECT 101.125 87.590 101.425 88.440 ;
        RECT 103.125 87.590 103.425 88.440 ;
        RECT 105.125 87.590 105.425 88.440 ;
        RECT 107.125 87.590 107.425 88.440 ;
        RECT 109.125 87.590 109.425 88.440 ;
        RECT 111.125 87.590 111.425 88.440 ;
        RECT 113.125 87.590 113.425 88.440 ;
        RECT 115.125 87.590 115.425 88.440 ;
        RECT 117.125 87.590 117.425 88.440 ;
        RECT 119.125 87.590 119.425 88.440 ;
        RECT 121.125 87.590 121.425 88.440 ;
        RECT 123.125 87.590 123.425 88.440 ;
        RECT 125.125 87.590 125.425 88.440 ;
        RECT 127.125 87.590 127.425 88.440 ;
        RECT 129.125 87.590 129.425 88.440 ;
        RECT 131.125 87.590 131.425 88.440 ;
        RECT 133.125 87.590 133.425 88.440 ;
        RECT 135.125 87.590 135.425 88.440 ;
        RECT 137.125 87.590 137.425 88.440 ;
        RECT 139.125 87.590 139.425 88.440 ;
        RECT 141.125 87.590 141.425 88.440 ;
        RECT 143.125 87.590 143.425 88.440 ;
        RECT 145.125 87.590 145.425 88.440 ;
        RECT 147.125 87.590 147.425 88.440 ;
        RECT 149.125 87.590 149.425 88.440 ;
        RECT 151.125 87.590 151.425 88.440 ;
        RECT 153.125 87.590 153.425 88.440 ;
        RECT 7.340 86.590 8.340 87.590 ;
        RECT 9.340 86.590 10.340 87.590 ;
        RECT 11.340 86.590 12.340 87.590 ;
        RECT 13.340 86.590 14.340 87.590 ;
        RECT 15.340 86.590 16.340 87.590 ;
        RECT 17.340 86.590 18.340 87.590 ;
        RECT 19.340 86.590 20.340 87.590 ;
        RECT 21.340 86.590 22.340 87.590 ;
        RECT 23.340 86.590 24.340 87.590 ;
        RECT 25.340 86.590 26.340 87.590 ;
        RECT 27.340 86.590 28.340 87.590 ;
        RECT 29.340 86.590 30.340 87.590 ;
        RECT 31.340 86.590 32.340 87.590 ;
        RECT 33.340 86.590 34.340 87.590 ;
        RECT 35.340 86.590 36.340 87.590 ;
        RECT 37.340 86.590 38.340 87.590 ;
        RECT 39.340 86.590 40.340 87.590 ;
        RECT 41.340 86.590 42.340 87.590 ;
        RECT 43.340 86.590 44.340 87.590 ;
        RECT 45.340 86.590 46.340 87.590 ;
        RECT 47.340 86.590 48.340 87.590 ;
        RECT 49.340 86.590 50.340 87.590 ;
        RECT 51.340 86.590 52.340 87.590 ;
        RECT 53.340 86.590 54.340 87.590 ;
        RECT 55.340 86.590 56.340 87.590 ;
        RECT 57.340 86.590 58.340 87.590 ;
        RECT 59.340 86.590 60.340 87.590 ;
        RECT 61.340 86.590 62.340 87.590 ;
        RECT 63.340 86.590 64.340 87.590 ;
        RECT 65.340 86.590 66.340 87.590 ;
        RECT 67.340 86.590 68.340 87.590 ;
        RECT 69.340 86.590 70.340 87.590 ;
        RECT 71.340 86.590 72.340 87.590 ;
        RECT 73.340 86.590 74.340 87.590 ;
        RECT 86.775 86.590 87.775 87.590 ;
        RECT 88.775 86.590 89.775 87.590 ;
        RECT 90.775 86.590 91.775 87.590 ;
        RECT 92.775 86.590 93.775 87.590 ;
        RECT 94.775 86.590 95.775 87.590 ;
        RECT 96.775 86.590 97.775 87.590 ;
        RECT 98.775 86.590 99.775 87.590 ;
        RECT 100.775 86.590 101.775 87.590 ;
        RECT 102.775 86.590 103.775 87.590 ;
        RECT 104.775 86.590 105.775 87.590 ;
        RECT 106.775 86.590 107.775 87.590 ;
        RECT 108.775 86.590 109.775 87.590 ;
        RECT 110.775 86.590 111.775 87.590 ;
        RECT 112.775 86.590 113.775 87.590 ;
        RECT 114.775 86.590 115.775 87.590 ;
        RECT 116.775 86.590 117.775 87.590 ;
        RECT 118.775 86.590 119.775 87.590 ;
        RECT 120.775 86.590 121.775 87.590 ;
        RECT 122.775 86.590 123.775 87.590 ;
        RECT 124.775 86.590 125.775 87.590 ;
        RECT 126.775 86.590 127.775 87.590 ;
        RECT 128.775 86.590 129.775 87.590 ;
        RECT 130.775 86.590 131.775 87.590 ;
        RECT 132.775 86.590 133.775 87.590 ;
        RECT 134.775 86.590 135.775 87.590 ;
        RECT 136.775 86.590 137.775 87.590 ;
        RECT 138.775 86.590 139.775 87.590 ;
        RECT 140.775 86.590 141.775 87.590 ;
        RECT 142.775 86.590 143.775 87.590 ;
        RECT 144.775 86.590 145.775 87.590 ;
        RECT 146.775 86.590 147.775 87.590 ;
        RECT 148.775 86.590 149.775 87.590 ;
        RECT 150.775 86.590 151.775 87.590 ;
        RECT 152.775 86.590 153.775 87.590 ;
        RECT 7.690 85.740 7.990 86.590 ;
        RECT 9.690 85.740 9.990 86.590 ;
        RECT 11.690 85.740 11.990 86.590 ;
        RECT 13.690 85.740 13.990 86.590 ;
        RECT 15.690 85.740 15.990 86.590 ;
        RECT 17.690 85.740 17.990 86.590 ;
        RECT 19.690 85.740 19.990 86.590 ;
        RECT 21.690 85.740 21.990 86.590 ;
        RECT 23.690 85.740 23.990 86.590 ;
        RECT 25.690 85.740 25.990 86.590 ;
        RECT 27.690 85.740 27.990 86.590 ;
        RECT 29.690 85.740 29.990 86.590 ;
        RECT 31.690 85.740 31.990 86.590 ;
        RECT 33.690 85.740 33.990 86.590 ;
        RECT 35.690 85.740 35.990 86.590 ;
        RECT 37.690 85.740 37.990 86.590 ;
        RECT 39.690 85.740 39.990 86.590 ;
        RECT 41.690 85.740 41.990 86.590 ;
        RECT 43.690 85.740 43.990 86.590 ;
        RECT 45.690 85.740 45.990 86.590 ;
        RECT 47.690 85.740 47.990 86.590 ;
        RECT 49.690 85.740 49.990 86.590 ;
        RECT 51.690 85.740 51.990 86.590 ;
        RECT 53.690 85.740 53.990 86.590 ;
        RECT 55.690 85.740 55.990 86.590 ;
        RECT 57.690 85.740 57.990 86.590 ;
        RECT 59.690 85.740 59.990 86.590 ;
        RECT 61.690 85.740 61.990 86.590 ;
        RECT 63.690 85.740 63.990 86.590 ;
        RECT 65.690 85.740 65.990 86.590 ;
        RECT 67.690 85.740 67.990 86.590 ;
        RECT 69.690 85.740 69.990 86.590 ;
        RECT 71.690 85.740 71.990 86.590 ;
        RECT 73.690 85.740 73.990 86.590 ;
        RECT 87.125 85.740 87.425 86.590 ;
        RECT 89.125 85.740 89.425 86.590 ;
        RECT 91.125 85.740 91.425 86.590 ;
        RECT 93.125 85.740 93.425 86.590 ;
        RECT 95.125 85.740 95.425 86.590 ;
        RECT 97.125 85.740 97.425 86.590 ;
        RECT 99.125 85.740 99.425 86.590 ;
        RECT 101.125 85.740 101.425 86.590 ;
        RECT 103.125 85.740 103.425 86.590 ;
        RECT 105.125 85.740 105.425 86.590 ;
        RECT 107.125 85.740 107.425 86.590 ;
        RECT 109.125 85.740 109.425 86.590 ;
        RECT 111.125 85.740 111.425 86.590 ;
        RECT 113.125 85.740 113.425 86.590 ;
        RECT 115.125 85.740 115.425 86.590 ;
        RECT 117.125 85.740 117.425 86.590 ;
        RECT 119.125 85.740 119.425 86.590 ;
        RECT 121.125 85.740 121.425 86.590 ;
        RECT 123.125 85.740 123.425 86.590 ;
        RECT 125.125 85.740 125.425 86.590 ;
        RECT 127.125 85.740 127.425 86.590 ;
        RECT 129.125 85.740 129.425 86.590 ;
        RECT 131.125 85.740 131.425 86.590 ;
        RECT 133.125 85.740 133.425 86.590 ;
        RECT 135.125 85.740 135.425 86.590 ;
        RECT 137.125 85.740 137.425 86.590 ;
        RECT 139.125 85.740 139.425 86.590 ;
        RECT 141.125 85.740 141.425 86.590 ;
        RECT 143.125 85.740 143.425 86.590 ;
        RECT 145.125 85.740 145.425 86.590 ;
        RECT 147.125 85.740 147.425 86.590 ;
        RECT 149.125 85.740 149.425 86.590 ;
        RECT 151.125 85.740 151.425 86.590 ;
        RECT 153.125 85.740 153.425 86.590 ;
        RECT 7.340 84.740 8.340 85.740 ;
        RECT 9.340 84.740 10.340 85.740 ;
        RECT 11.340 84.740 12.340 85.740 ;
        RECT 13.340 84.740 14.340 85.740 ;
        RECT 15.340 84.740 16.340 85.740 ;
        RECT 17.340 84.740 18.340 85.740 ;
        RECT 19.340 84.740 20.340 85.740 ;
        RECT 21.340 84.740 22.340 85.740 ;
        RECT 23.340 84.740 24.340 85.740 ;
        RECT 25.340 84.740 26.340 85.740 ;
        RECT 27.340 84.740 28.340 85.740 ;
        RECT 29.340 84.740 30.340 85.740 ;
        RECT 31.340 84.740 32.340 85.740 ;
        RECT 33.340 84.740 34.340 85.740 ;
        RECT 35.340 84.740 36.340 85.740 ;
        RECT 37.340 84.740 38.340 85.740 ;
        RECT 39.340 84.740 40.340 85.740 ;
        RECT 41.340 84.740 42.340 85.740 ;
        RECT 43.340 84.740 44.340 85.740 ;
        RECT 45.340 84.740 46.340 85.740 ;
        RECT 47.340 84.740 48.340 85.740 ;
        RECT 49.340 84.740 50.340 85.740 ;
        RECT 51.340 84.740 52.340 85.740 ;
        RECT 53.340 84.740 54.340 85.740 ;
        RECT 55.340 84.740 56.340 85.740 ;
        RECT 57.340 84.740 58.340 85.740 ;
        RECT 59.340 84.740 60.340 85.740 ;
        RECT 61.340 84.740 62.340 85.740 ;
        RECT 63.340 84.740 64.340 85.740 ;
        RECT 65.340 84.740 66.340 85.740 ;
        RECT 67.340 84.740 68.340 85.740 ;
        RECT 69.340 84.740 70.340 85.740 ;
        RECT 71.340 84.740 72.340 85.740 ;
        RECT 73.340 84.740 74.340 85.740 ;
        RECT 86.775 84.740 87.775 85.740 ;
        RECT 88.775 84.740 89.775 85.740 ;
        RECT 90.775 84.740 91.775 85.740 ;
        RECT 92.775 84.740 93.775 85.740 ;
        RECT 94.775 84.740 95.775 85.740 ;
        RECT 96.775 84.740 97.775 85.740 ;
        RECT 98.775 84.740 99.775 85.740 ;
        RECT 100.775 84.740 101.775 85.740 ;
        RECT 102.775 84.740 103.775 85.740 ;
        RECT 104.775 84.740 105.775 85.740 ;
        RECT 106.775 84.740 107.775 85.740 ;
        RECT 108.775 84.740 109.775 85.740 ;
        RECT 110.775 84.740 111.775 85.740 ;
        RECT 112.775 84.740 113.775 85.740 ;
        RECT 114.775 84.740 115.775 85.740 ;
        RECT 116.775 84.740 117.775 85.740 ;
        RECT 118.775 84.740 119.775 85.740 ;
        RECT 120.775 84.740 121.775 85.740 ;
        RECT 122.775 84.740 123.775 85.740 ;
        RECT 124.775 84.740 125.775 85.740 ;
        RECT 126.775 84.740 127.775 85.740 ;
        RECT 128.775 84.740 129.775 85.740 ;
        RECT 130.775 84.740 131.775 85.740 ;
        RECT 132.775 84.740 133.775 85.740 ;
        RECT 134.775 84.740 135.775 85.740 ;
        RECT 136.775 84.740 137.775 85.740 ;
        RECT 138.775 84.740 139.775 85.740 ;
        RECT 140.775 84.740 141.775 85.740 ;
        RECT 142.775 84.740 143.775 85.740 ;
        RECT 144.775 84.740 145.775 85.740 ;
        RECT 146.775 84.740 147.775 85.740 ;
        RECT 148.775 84.740 149.775 85.740 ;
        RECT 150.775 84.740 151.775 85.740 ;
        RECT 152.775 84.740 153.775 85.740 ;
        RECT 7.690 83.890 7.990 84.740 ;
        RECT 9.690 83.890 9.990 84.740 ;
        RECT 11.690 83.890 11.990 84.740 ;
        RECT 13.690 83.890 13.990 84.740 ;
        RECT 15.690 83.890 15.990 84.740 ;
        RECT 17.690 83.890 17.990 84.740 ;
        RECT 19.690 83.890 19.990 84.740 ;
        RECT 21.690 83.890 21.990 84.740 ;
        RECT 23.690 83.890 23.990 84.740 ;
        RECT 25.690 83.890 25.990 84.740 ;
        RECT 27.690 83.890 27.990 84.740 ;
        RECT 29.690 83.890 29.990 84.740 ;
        RECT 31.690 83.890 31.990 84.740 ;
        RECT 33.690 83.890 33.990 84.740 ;
        RECT 35.690 83.890 35.990 84.740 ;
        RECT 37.690 83.890 37.990 84.740 ;
        RECT 39.690 83.890 39.990 84.740 ;
        RECT 41.690 83.890 41.990 84.740 ;
        RECT 43.690 83.890 43.990 84.740 ;
        RECT 45.690 83.890 45.990 84.740 ;
        RECT 47.690 83.890 47.990 84.740 ;
        RECT 49.690 83.890 49.990 84.740 ;
        RECT 51.690 83.890 51.990 84.740 ;
        RECT 53.690 83.890 53.990 84.740 ;
        RECT 55.690 83.890 55.990 84.740 ;
        RECT 57.690 83.890 57.990 84.740 ;
        RECT 59.690 83.890 59.990 84.740 ;
        RECT 61.690 83.890 61.990 84.740 ;
        RECT 63.690 83.890 63.990 84.740 ;
        RECT 65.690 83.890 65.990 84.740 ;
        RECT 67.690 83.890 67.990 84.740 ;
        RECT 69.690 83.890 69.990 84.740 ;
        RECT 71.690 83.890 71.990 84.740 ;
        RECT 73.690 83.890 73.990 84.740 ;
        RECT 87.125 83.890 87.425 84.740 ;
        RECT 89.125 83.890 89.425 84.740 ;
        RECT 91.125 83.890 91.425 84.740 ;
        RECT 93.125 83.890 93.425 84.740 ;
        RECT 95.125 83.890 95.425 84.740 ;
        RECT 97.125 83.890 97.425 84.740 ;
        RECT 99.125 83.890 99.425 84.740 ;
        RECT 101.125 83.890 101.425 84.740 ;
        RECT 103.125 83.890 103.425 84.740 ;
        RECT 105.125 83.890 105.425 84.740 ;
        RECT 107.125 83.890 107.425 84.740 ;
        RECT 109.125 83.890 109.425 84.740 ;
        RECT 111.125 83.890 111.425 84.740 ;
        RECT 113.125 83.890 113.425 84.740 ;
        RECT 115.125 83.890 115.425 84.740 ;
        RECT 117.125 83.890 117.425 84.740 ;
        RECT 119.125 83.890 119.425 84.740 ;
        RECT 121.125 83.890 121.425 84.740 ;
        RECT 123.125 83.890 123.425 84.740 ;
        RECT 125.125 83.890 125.425 84.740 ;
        RECT 127.125 83.890 127.425 84.740 ;
        RECT 129.125 83.890 129.425 84.740 ;
        RECT 131.125 83.890 131.425 84.740 ;
        RECT 133.125 83.890 133.425 84.740 ;
        RECT 135.125 83.890 135.425 84.740 ;
        RECT 137.125 83.890 137.425 84.740 ;
        RECT 139.125 83.890 139.425 84.740 ;
        RECT 141.125 83.890 141.425 84.740 ;
        RECT 143.125 83.890 143.425 84.740 ;
        RECT 145.125 83.890 145.425 84.740 ;
        RECT 147.125 83.890 147.425 84.740 ;
        RECT 149.125 83.890 149.425 84.740 ;
        RECT 151.125 83.890 151.425 84.740 ;
        RECT 153.125 83.890 153.425 84.740 ;
        RECT 7.340 82.890 8.340 83.890 ;
        RECT 9.340 82.890 10.340 83.890 ;
        RECT 11.340 82.890 12.340 83.890 ;
        RECT 13.340 82.890 14.340 83.890 ;
        RECT 15.340 82.890 16.340 83.890 ;
        RECT 17.340 82.890 18.340 83.890 ;
        RECT 19.340 82.890 20.340 83.890 ;
        RECT 21.340 82.890 22.340 83.890 ;
        RECT 23.340 82.890 24.340 83.890 ;
        RECT 25.340 82.890 26.340 83.890 ;
        RECT 27.340 82.890 28.340 83.890 ;
        RECT 29.340 82.890 30.340 83.890 ;
        RECT 31.340 82.890 32.340 83.890 ;
        RECT 33.340 82.890 34.340 83.890 ;
        RECT 35.340 82.890 36.340 83.890 ;
        RECT 37.340 82.890 38.340 83.890 ;
        RECT 39.340 82.890 40.340 83.890 ;
        RECT 41.340 82.890 42.340 83.890 ;
        RECT 43.340 82.890 44.340 83.890 ;
        RECT 45.340 82.890 46.340 83.890 ;
        RECT 47.340 82.890 48.340 83.890 ;
        RECT 49.340 82.890 50.340 83.890 ;
        RECT 51.340 82.890 52.340 83.890 ;
        RECT 53.340 82.890 54.340 83.890 ;
        RECT 55.340 82.890 56.340 83.890 ;
        RECT 57.340 82.890 58.340 83.890 ;
        RECT 59.340 82.890 60.340 83.890 ;
        RECT 61.340 82.890 62.340 83.890 ;
        RECT 63.340 82.890 64.340 83.890 ;
        RECT 65.340 82.890 66.340 83.890 ;
        RECT 67.340 82.890 68.340 83.890 ;
        RECT 69.340 82.890 70.340 83.890 ;
        RECT 71.340 82.890 72.340 83.890 ;
        RECT 73.340 82.890 74.340 83.890 ;
        RECT 86.775 82.890 87.775 83.890 ;
        RECT 88.775 82.890 89.775 83.890 ;
        RECT 90.775 82.890 91.775 83.890 ;
        RECT 92.775 82.890 93.775 83.890 ;
        RECT 94.775 82.890 95.775 83.890 ;
        RECT 96.775 82.890 97.775 83.890 ;
        RECT 98.775 82.890 99.775 83.890 ;
        RECT 100.775 82.890 101.775 83.890 ;
        RECT 102.775 82.890 103.775 83.890 ;
        RECT 104.775 82.890 105.775 83.890 ;
        RECT 106.775 82.890 107.775 83.890 ;
        RECT 108.775 82.890 109.775 83.890 ;
        RECT 110.775 82.890 111.775 83.890 ;
        RECT 112.775 82.890 113.775 83.890 ;
        RECT 114.775 82.890 115.775 83.890 ;
        RECT 116.775 82.890 117.775 83.890 ;
        RECT 118.775 82.890 119.775 83.890 ;
        RECT 120.775 82.890 121.775 83.890 ;
        RECT 122.775 82.890 123.775 83.890 ;
        RECT 124.775 82.890 125.775 83.890 ;
        RECT 126.775 82.890 127.775 83.890 ;
        RECT 128.775 82.890 129.775 83.890 ;
        RECT 130.775 82.890 131.775 83.890 ;
        RECT 132.775 82.890 133.775 83.890 ;
        RECT 134.775 82.890 135.775 83.890 ;
        RECT 136.775 82.890 137.775 83.890 ;
        RECT 138.775 82.890 139.775 83.890 ;
        RECT 140.775 82.890 141.775 83.890 ;
        RECT 142.775 82.890 143.775 83.890 ;
        RECT 144.775 82.890 145.775 83.890 ;
        RECT 146.775 82.890 147.775 83.890 ;
        RECT 148.775 82.890 149.775 83.890 ;
        RECT 150.775 82.890 151.775 83.890 ;
        RECT 152.775 82.890 153.775 83.890 ;
        RECT 7.690 82.040 7.990 82.890 ;
        RECT 9.690 82.040 9.990 82.890 ;
        RECT 11.690 82.040 11.990 82.890 ;
        RECT 13.690 82.040 13.990 82.890 ;
        RECT 15.690 82.040 15.990 82.890 ;
        RECT 17.690 82.040 17.990 82.890 ;
        RECT 19.690 82.040 19.990 82.890 ;
        RECT 21.690 82.040 21.990 82.890 ;
        RECT 23.690 82.040 23.990 82.890 ;
        RECT 25.690 82.040 25.990 82.890 ;
        RECT 27.690 82.040 27.990 82.890 ;
        RECT 29.690 82.040 29.990 82.890 ;
        RECT 31.690 82.040 31.990 82.890 ;
        RECT 33.690 82.040 33.990 82.890 ;
        RECT 35.690 82.040 35.990 82.890 ;
        RECT 37.690 82.040 37.990 82.890 ;
        RECT 39.690 82.040 39.990 82.890 ;
        RECT 41.690 82.040 41.990 82.890 ;
        RECT 43.690 82.040 43.990 82.890 ;
        RECT 45.690 82.040 45.990 82.890 ;
        RECT 47.690 82.040 47.990 82.890 ;
        RECT 49.690 82.040 49.990 82.890 ;
        RECT 51.690 82.040 51.990 82.890 ;
        RECT 53.690 82.040 53.990 82.890 ;
        RECT 55.690 82.040 55.990 82.890 ;
        RECT 57.690 82.040 57.990 82.890 ;
        RECT 59.690 82.040 59.990 82.890 ;
        RECT 61.690 82.040 61.990 82.890 ;
        RECT 63.690 82.040 63.990 82.890 ;
        RECT 65.690 82.040 65.990 82.890 ;
        RECT 67.690 82.040 67.990 82.890 ;
        RECT 69.690 82.040 69.990 82.890 ;
        RECT 71.690 82.040 71.990 82.890 ;
        RECT 73.690 82.040 73.990 82.890 ;
        RECT 87.125 82.040 87.425 82.890 ;
        RECT 89.125 82.040 89.425 82.890 ;
        RECT 91.125 82.040 91.425 82.890 ;
        RECT 93.125 82.040 93.425 82.890 ;
        RECT 95.125 82.040 95.425 82.890 ;
        RECT 97.125 82.040 97.425 82.890 ;
        RECT 99.125 82.040 99.425 82.890 ;
        RECT 101.125 82.040 101.425 82.890 ;
        RECT 103.125 82.040 103.425 82.890 ;
        RECT 105.125 82.040 105.425 82.890 ;
        RECT 107.125 82.040 107.425 82.890 ;
        RECT 109.125 82.040 109.425 82.890 ;
        RECT 111.125 82.040 111.425 82.890 ;
        RECT 113.125 82.040 113.425 82.890 ;
        RECT 115.125 82.040 115.425 82.890 ;
        RECT 117.125 82.040 117.425 82.890 ;
        RECT 119.125 82.040 119.425 82.890 ;
        RECT 121.125 82.040 121.425 82.890 ;
        RECT 123.125 82.040 123.425 82.890 ;
        RECT 125.125 82.040 125.425 82.890 ;
        RECT 127.125 82.040 127.425 82.890 ;
        RECT 129.125 82.040 129.425 82.890 ;
        RECT 131.125 82.040 131.425 82.890 ;
        RECT 133.125 82.040 133.425 82.890 ;
        RECT 135.125 82.040 135.425 82.890 ;
        RECT 137.125 82.040 137.425 82.890 ;
        RECT 139.125 82.040 139.425 82.890 ;
        RECT 141.125 82.040 141.425 82.890 ;
        RECT 143.125 82.040 143.425 82.890 ;
        RECT 145.125 82.040 145.425 82.890 ;
        RECT 147.125 82.040 147.425 82.890 ;
        RECT 149.125 82.040 149.425 82.890 ;
        RECT 151.125 82.040 151.425 82.890 ;
        RECT 153.125 82.040 153.425 82.890 ;
        RECT 7.340 81.040 8.340 82.040 ;
        RECT 9.340 81.040 10.340 82.040 ;
        RECT 11.340 81.040 12.340 82.040 ;
        RECT 13.340 81.040 14.340 82.040 ;
        RECT 15.340 81.040 16.340 82.040 ;
        RECT 17.340 81.040 18.340 82.040 ;
        RECT 19.340 81.040 20.340 82.040 ;
        RECT 21.340 81.040 22.340 82.040 ;
        RECT 23.340 81.040 24.340 82.040 ;
        RECT 25.340 81.040 26.340 82.040 ;
        RECT 27.340 81.040 28.340 82.040 ;
        RECT 29.340 81.040 30.340 82.040 ;
        RECT 31.340 81.040 32.340 82.040 ;
        RECT 33.340 81.040 34.340 82.040 ;
        RECT 35.340 81.040 36.340 82.040 ;
        RECT 37.340 81.040 38.340 82.040 ;
        RECT 39.340 81.040 40.340 82.040 ;
        RECT 41.340 81.040 42.340 82.040 ;
        RECT 43.340 81.040 44.340 82.040 ;
        RECT 45.340 81.040 46.340 82.040 ;
        RECT 47.340 81.040 48.340 82.040 ;
        RECT 49.340 81.040 50.340 82.040 ;
        RECT 51.340 81.040 52.340 82.040 ;
        RECT 53.340 81.040 54.340 82.040 ;
        RECT 55.340 81.040 56.340 82.040 ;
        RECT 57.340 81.040 58.340 82.040 ;
        RECT 59.340 81.040 60.340 82.040 ;
        RECT 61.340 81.040 62.340 82.040 ;
        RECT 63.340 81.040 64.340 82.040 ;
        RECT 65.340 81.040 66.340 82.040 ;
        RECT 67.340 81.040 68.340 82.040 ;
        RECT 69.340 81.040 70.340 82.040 ;
        RECT 71.340 81.040 72.340 82.040 ;
        RECT 73.340 81.040 74.340 82.040 ;
        RECT 86.775 81.040 87.775 82.040 ;
        RECT 88.775 81.040 89.775 82.040 ;
        RECT 90.775 81.040 91.775 82.040 ;
        RECT 92.775 81.040 93.775 82.040 ;
        RECT 94.775 81.040 95.775 82.040 ;
        RECT 96.775 81.040 97.775 82.040 ;
        RECT 98.775 81.040 99.775 82.040 ;
        RECT 100.775 81.040 101.775 82.040 ;
        RECT 102.775 81.040 103.775 82.040 ;
        RECT 104.775 81.040 105.775 82.040 ;
        RECT 106.775 81.040 107.775 82.040 ;
        RECT 108.775 81.040 109.775 82.040 ;
        RECT 110.775 81.040 111.775 82.040 ;
        RECT 112.775 81.040 113.775 82.040 ;
        RECT 114.775 81.040 115.775 82.040 ;
        RECT 116.775 81.040 117.775 82.040 ;
        RECT 118.775 81.040 119.775 82.040 ;
        RECT 120.775 81.040 121.775 82.040 ;
        RECT 122.775 81.040 123.775 82.040 ;
        RECT 124.775 81.040 125.775 82.040 ;
        RECT 126.775 81.040 127.775 82.040 ;
        RECT 128.775 81.040 129.775 82.040 ;
        RECT 130.775 81.040 131.775 82.040 ;
        RECT 132.775 81.040 133.775 82.040 ;
        RECT 134.775 81.040 135.775 82.040 ;
        RECT 136.775 81.040 137.775 82.040 ;
        RECT 138.775 81.040 139.775 82.040 ;
        RECT 140.775 81.040 141.775 82.040 ;
        RECT 142.775 81.040 143.775 82.040 ;
        RECT 144.775 81.040 145.775 82.040 ;
        RECT 146.775 81.040 147.775 82.040 ;
        RECT 148.775 81.040 149.775 82.040 ;
        RECT 150.775 81.040 151.775 82.040 ;
        RECT 152.775 81.040 153.775 82.040 ;
        RECT 7.690 80.190 7.990 81.040 ;
        RECT 9.690 80.190 9.990 81.040 ;
        RECT 11.690 80.190 11.990 81.040 ;
        RECT 13.690 80.190 13.990 81.040 ;
        RECT 15.690 80.190 15.990 81.040 ;
        RECT 17.690 80.190 17.990 81.040 ;
        RECT 19.690 80.190 19.990 81.040 ;
        RECT 21.690 80.190 21.990 81.040 ;
        RECT 23.690 80.190 23.990 81.040 ;
        RECT 25.690 80.190 25.990 81.040 ;
        RECT 27.690 80.190 27.990 81.040 ;
        RECT 29.690 80.190 29.990 81.040 ;
        RECT 31.690 80.190 31.990 81.040 ;
        RECT 33.690 80.190 33.990 81.040 ;
        RECT 35.690 80.190 35.990 81.040 ;
        RECT 37.690 80.190 37.990 81.040 ;
        RECT 39.690 80.190 39.990 81.040 ;
        RECT 41.690 80.190 41.990 81.040 ;
        RECT 43.690 80.190 43.990 81.040 ;
        RECT 45.690 80.190 45.990 81.040 ;
        RECT 47.690 80.190 47.990 81.040 ;
        RECT 49.690 80.190 49.990 81.040 ;
        RECT 51.690 80.190 51.990 81.040 ;
        RECT 53.690 80.190 53.990 81.040 ;
        RECT 55.690 80.190 55.990 81.040 ;
        RECT 57.690 80.190 57.990 81.040 ;
        RECT 59.690 80.190 59.990 81.040 ;
        RECT 61.690 80.190 61.990 81.040 ;
        RECT 63.690 80.190 63.990 81.040 ;
        RECT 65.690 80.190 65.990 81.040 ;
        RECT 67.690 80.190 67.990 81.040 ;
        RECT 69.690 80.190 69.990 81.040 ;
        RECT 71.690 80.190 71.990 81.040 ;
        RECT 73.690 80.190 73.990 81.040 ;
        RECT 87.125 80.190 87.425 81.040 ;
        RECT 89.125 80.190 89.425 81.040 ;
        RECT 91.125 80.190 91.425 81.040 ;
        RECT 93.125 80.190 93.425 81.040 ;
        RECT 95.125 80.190 95.425 81.040 ;
        RECT 97.125 80.190 97.425 81.040 ;
        RECT 99.125 80.190 99.425 81.040 ;
        RECT 101.125 80.190 101.425 81.040 ;
        RECT 103.125 80.190 103.425 81.040 ;
        RECT 105.125 80.190 105.425 81.040 ;
        RECT 107.125 80.190 107.425 81.040 ;
        RECT 109.125 80.190 109.425 81.040 ;
        RECT 111.125 80.190 111.425 81.040 ;
        RECT 113.125 80.190 113.425 81.040 ;
        RECT 115.125 80.190 115.425 81.040 ;
        RECT 117.125 80.190 117.425 81.040 ;
        RECT 119.125 80.190 119.425 81.040 ;
        RECT 121.125 80.190 121.425 81.040 ;
        RECT 123.125 80.190 123.425 81.040 ;
        RECT 125.125 80.190 125.425 81.040 ;
        RECT 127.125 80.190 127.425 81.040 ;
        RECT 129.125 80.190 129.425 81.040 ;
        RECT 131.125 80.190 131.425 81.040 ;
        RECT 133.125 80.190 133.425 81.040 ;
        RECT 135.125 80.190 135.425 81.040 ;
        RECT 137.125 80.190 137.425 81.040 ;
        RECT 139.125 80.190 139.425 81.040 ;
        RECT 141.125 80.190 141.425 81.040 ;
        RECT 143.125 80.190 143.425 81.040 ;
        RECT 145.125 80.190 145.425 81.040 ;
        RECT 147.125 80.190 147.425 81.040 ;
        RECT 149.125 80.190 149.425 81.040 ;
        RECT 151.125 80.190 151.425 81.040 ;
        RECT 153.125 80.190 153.425 81.040 ;
        RECT 7.340 79.190 8.340 80.190 ;
        RECT 9.340 79.190 10.340 80.190 ;
        RECT 11.340 79.190 12.340 80.190 ;
        RECT 13.340 79.190 14.340 80.190 ;
        RECT 15.340 79.190 16.340 80.190 ;
        RECT 17.340 79.190 18.340 80.190 ;
        RECT 19.340 79.190 20.340 80.190 ;
        RECT 21.340 79.190 22.340 80.190 ;
        RECT 23.340 79.190 24.340 80.190 ;
        RECT 25.340 79.190 26.340 80.190 ;
        RECT 27.340 79.190 28.340 80.190 ;
        RECT 29.340 79.190 30.340 80.190 ;
        RECT 31.340 79.190 32.340 80.190 ;
        RECT 33.340 79.190 34.340 80.190 ;
        RECT 35.340 79.190 36.340 80.190 ;
        RECT 37.340 79.190 38.340 80.190 ;
        RECT 39.340 79.190 40.340 80.190 ;
        RECT 41.340 79.190 42.340 80.190 ;
        RECT 43.340 79.190 44.340 80.190 ;
        RECT 45.340 79.190 46.340 80.190 ;
        RECT 47.340 79.190 48.340 80.190 ;
        RECT 49.340 79.190 50.340 80.190 ;
        RECT 51.340 79.190 52.340 80.190 ;
        RECT 53.340 79.190 54.340 80.190 ;
        RECT 55.340 79.190 56.340 80.190 ;
        RECT 57.340 79.190 58.340 80.190 ;
        RECT 59.340 79.190 60.340 80.190 ;
        RECT 61.340 79.190 62.340 80.190 ;
        RECT 63.340 79.190 64.340 80.190 ;
        RECT 65.340 79.190 66.340 80.190 ;
        RECT 67.340 79.190 68.340 80.190 ;
        RECT 69.340 79.190 70.340 80.190 ;
        RECT 71.340 79.190 72.340 80.190 ;
        RECT 73.340 79.190 74.340 80.190 ;
        RECT 86.775 79.190 87.775 80.190 ;
        RECT 88.775 79.190 89.775 80.190 ;
        RECT 90.775 79.190 91.775 80.190 ;
        RECT 92.775 79.190 93.775 80.190 ;
        RECT 94.775 79.190 95.775 80.190 ;
        RECT 96.775 79.190 97.775 80.190 ;
        RECT 98.775 79.190 99.775 80.190 ;
        RECT 100.775 79.190 101.775 80.190 ;
        RECT 102.775 79.190 103.775 80.190 ;
        RECT 104.775 79.190 105.775 80.190 ;
        RECT 106.775 79.190 107.775 80.190 ;
        RECT 108.775 79.190 109.775 80.190 ;
        RECT 110.775 79.190 111.775 80.190 ;
        RECT 112.775 79.190 113.775 80.190 ;
        RECT 114.775 79.190 115.775 80.190 ;
        RECT 116.775 79.190 117.775 80.190 ;
        RECT 118.775 79.190 119.775 80.190 ;
        RECT 120.775 79.190 121.775 80.190 ;
        RECT 122.775 79.190 123.775 80.190 ;
        RECT 124.775 79.190 125.775 80.190 ;
        RECT 126.775 79.190 127.775 80.190 ;
        RECT 128.775 79.190 129.775 80.190 ;
        RECT 130.775 79.190 131.775 80.190 ;
        RECT 132.775 79.190 133.775 80.190 ;
        RECT 134.775 79.190 135.775 80.190 ;
        RECT 136.775 79.190 137.775 80.190 ;
        RECT 138.775 79.190 139.775 80.190 ;
        RECT 140.775 79.190 141.775 80.190 ;
        RECT 142.775 79.190 143.775 80.190 ;
        RECT 144.775 79.190 145.775 80.190 ;
        RECT 146.775 79.190 147.775 80.190 ;
        RECT 148.775 79.190 149.775 80.190 ;
        RECT 150.775 79.190 151.775 80.190 ;
        RECT 152.775 79.190 153.775 80.190 ;
        RECT 7.690 78.340 7.990 79.190 ;
        RECT 9.690 78.340 9.990 79.190 ;
        RECT 11.690 78.340 11.990 79.190 ;
        RECT 13.690 78.340 13.990 79.190 ;
        RECT 15.690 78.340 15.990 79.190 ;
        RECT 17.690 78.340 17.990 79.190 ;
        RECT 19.690 78.340 19.990 79.190 ;
        RECT 21.690 78.340 21.990 79.190 ;
        RECT 23.690 78.340 23.990 79.190 ;
        RECT 25.690 78.340 25.990 79.190 ;
        RECT 27.690 78.340 27.990 79.190 ;
        RECT 29.690 78.340 29.990 79.190 ;
        RECT 31.690 78.340 31.990 79.190 ;
        RECT 33.690 78.340 33.990 79.190 ;
        RECT 35.690 78.340 35.990 79.190 ;
        RECT 37.690 78.340 37.990 79.190 ;
        RECT 39.690 78.340 39.990 79.190 ;
        RECT 41.690 78.340 41.990 79.190 ;
        RECT 43.690 78.340 43.990 79.190 ;
        RECT 45.690 78.340 45.990 79.190 ;
        RECT 47.690 78.340 47.990 79.190 ;
        RECT 49.690 78.340 49.990 79.190 ;
        RECT 51.690 78.340 51.990 79.190 ;
        RECT 53.690 78.340 53.990 79.190 ;
        RECT 55.690 78.340 55.990 79.190 ;
        RECT 57.690 78.340 57.990 79.190 ;
        RECT 59.690 78.340 59.990 79.190 ;
        RECT 61.690 78.340 61.990 79.190 ;
        RECT 63.690 78.340 63.990 79.190 ;
        RECT 65.690 78.340 65.990 79.190 ;
        RECT 67.690 78.340 67.990 79.190 ;
        RECT 69.690 78.340 69.990 79.190 ;
        RECT 71.690 78.340 71.990 79.190 ;
        RECT 73.690 78.340 73.990 79.190 ;
        RECT 87.125 78.340 87.425 79.190 ;
        RECT 89.125 78.340 89.425 79.190 ;
        RECT 91.125 78.340 91.425 79.190 ;
        RECT 93.125 78.340 93.425 79.190 ;
        RECT 95.125 78.340 95.425 79.190 ;
        RECT 97.125 78.340 97.425 79.190 ;
        RECT 99.125 78.340 99.425 79.190 ;
        RECT 101.125 78.340 101.425 79.190 ;
        RECT 103.125 78.340 103.425 79.190 ;
        RECT 105.125 78.340 105.425 79.190 ;
        RECT 107.125 78.340 107.425 79.190 ;
        RECT 109.125 78.340 109.425 79.190 ;
        RECT 111.125 78.340 111.425 79.190 ;
        RECT 113.125 78.340 113.425 79.190 ;
        RECT 115.125 78.340 115.425 79.190 ;
        RECT 117.125 78.340 117.425 79.190 ;
        RECT 119.125 78.340 119.425 79.190 ;
        RECT 121.125 78.340 121.425 79.190 ;
        RECT 123.125 78.340 123.425 79.190 ;
        RECT 125.125 78.340 125.425 79.190 ;
        RECT 127.125 78.340 127.425 79.190 ;
        RECT 129.125 78.340 129.425 79.190 ;
        RECT 131.125 78.340 131.425 79.190 ;
        RECT 133.125 78.340 133.425 79.190 ;
        RECT 135.125 78.340 135.425 79.190 ;
        RECT 137.125 78.340 137.425 79.190 ;
        RECT 139.125 78.340 139.425 79.190 ;
        RECT 141.125 78.340 141.425 79.190 ;
        RECT 143.125 78.340 143.425 79.190 ;
        RECT 145.125 78.340 145.425 79.190 ;
        RECT 147.125 78.340 147.425 79.190 ;
        RECT 149.125 78.340 149.425 79.190 ;
        RECT 151.125 78.340 151.425 79.190 ;
        RECT 153.125 78.340 153.425 79.190 ;
        RECT 7.340 77.340 8.340 78.340 ;
        RECT 9.340 77.340 10.340 78.340 ;
        RECT 11.340 77.340 12.340 78.340 ;
        RECT 13.340 77.340 14.340 78.340 ;
        RECT 15.340 77.340 16.340 78.340 ;
        RECT 17.340 77.340 18.340 78.340 ;
        RECT 19.340 77.340 20.340 78.340 ;
        RECT 21.340 77.340 22.340 78.340 ;
        RECT 23.340 77.340 24.340 78.340 ;
        RECT 25.340 77.340 26.340 78.340 ;
        RECT 27.340 77.340 28.340 78.340 ;
        RECT 29.340 77.340 30.340 78.340 ;
        RECT 31.340 77.340 32.340 78.340 ;
        RECT 33.340 77.340 34.340 78.340 ;
        RECT 35.340 77.340 36.340 78.340 ;
        RECT 37.340 77.340 38.340 78.340 ;
        RECT 39.340 77.340 40.340 78.340 ;
        RECT 41.340 77.340 42.340 78.340 ;
        RECT 43.340 77.340 44.340 78.340 ;
        RECT 45.340 77.340 46.340 78.340 ;
        RECT 47.340 77.340 48.340 78.340 ;
        RECT 49.340 77.340 50.340 78.340 ;
        RECT 51.340 77.340 52.340 78.340 ;
        RECT 53.340 77.340 54.340 78.340 ;
        RECT 55.340 77.340 56.340 78.340 ;
        RECT 57.340 77.340 58.340 78.340 ;
        RECT 59.340 77.340 60.340 78.340 ;
        RECT 61.340 77.340 62.340 78.340 ;
        RECT 63.340 77.340 64.340 78.340 ;
        RECT 65.340 77.340 66.340 78.340 ;
        RECT 67.340 77.340 68.340 78.340 ;
        RECT 69.340 77.340 70.340 78.340 ;
        RECT 71.340 77.340 72.340 78.340 ;
        RECT 73.340 77.340 74.340 78.340 ;
        RECT 86.775 77.340 87.775 78.340 ;
        RECT 88.775 77.340 89.775 78.340 ;
        RECT 90.775 77.340 91.775 78.340 ;
        RECT 92.775 77.340 93.775 78.340 ;
        RECT 94.775 77.340 95.775 78.340 ;
        RECT 96.775 77.340 97.775 78.340 ;
        RECT 98.775 77.340 99.775 78.340 ;
        RECT 100.775 77.340 101.775 78.340 ;
        RECT 102.775 77.340 103.775 78.340 ;
        RECT 104.775 77.340 105.775 78.340 ;
        RECT 106.775 77.340 107.775 78.340 ;
        RECT 108.775 77.340 109.775 78.340 ;
        RECT 110.775 77.340 111.775 78.340 ;
        RECT 112.775 77.340 113.775 78.340 ;
        RECT 114.775 77.340 115.775 78.340 ;
        RECT 116.775 77.340 117.775 78.340 ;
        RECT 118.775 77.340 119.775 78.340 ;
        RECT 120.775 77.340 121.775 78.340 ;
        RECT 122.775 77.340 123.775 78.340 ;
        RECT 124.775 77.340 125.775 78.340 ;
        RECT 126.775 77.340 127.775 78.340 ;
        RECT 128.775 77.340 129.775 78.340 ;
        RECT 130.775 77.340 131.775 78.340 ;
        RECT 132.775 77.340 133.775 78.340 ;
        RECT 134.775 77.340 135.775 78.340 ;
        RECT 136.775 77.340 137.775 78.340 ;
        RECT 138.775 77.340 139.775 78.340 ;
        RECT 140.775 77.340 141.775 78.340 ;
        RECT 142.775 77.340 143.775 78.340 ;
        RECT 144.775 77.340 145.775 78.340 ;
        RECT 146.775 77.340 147.775 78.340 ;
        RECT 148.775 77.340 149.775 78.340 ;
        RECT 150.775 77.340 151.775 78.340 ;
        RECT 152.775 77.340 153.775 78.340 ;
        RECT 7.690 76.490 7.990 77.340 ;
        RECT 9.690 76.490 9.990 77.340 ;
        RECT 11.690 76.490 11.990 77.340 ;
        RECT 13.690 76.490 13.990 77.340 ;
        RECT 15.690 76.490 15.990 77.340 ;
        RECT 17.690 76.490 17.990 77.340 ;
        RECT 19.690 76.490 19.990 77.340 ;
        RECT 21.690 76.490 21.990 77.340 ;
        RECT 23.690 76.490 23.990 77.340 ;
        RECT 25.690 76.490 25.990 77.340 ;
        RECT 27.690 76.490 27.990 77.340 ;
        RECT 29.690 76.490 29.990 77.340 ;
        RECT 31.690 76.490 31.990 77.340 ;
        RECT 33.690 76.490 33.990 77.340 ;
        RECT 35.690 76.490 35.990 77.340 ;
        RECT 37.690 76.490 37.990 77.340 ;
        RECT 39.690 76.490 39.990 77.340 ;
        RECT 41.690 76.490 41.990 77.340 ;
        RECT 43.690 76.490 43.990 77.340 ;
        RECT 45.690 76.490 45.990 77.340 ;
        RECT 47.690 76.490 47.990 77.340 ;
        RECT 49.690 76.490 49.990 77.340 ;
        RECT 51.690 76.490 51.990 77.340 ;
        RECT 53.690 76.490 53.990 77.340 ;
        RECT 55.690 76.490 55.990 77.340 ;
        RECT 57.690 76.490 57.990 77.340 ;
        RECT 59.690 76.490 59.990 77.340 ;
        RECT 61.690 76.490 61.990 77.340 ;
        RECT 63.690 76.490 63.990 77.340 ;
        RECT 65.690 76.490 65.990 77.340 ;
        RECT 67.690 76.490 67.990 77.340 ;
        RECT 69.690 76.490 69.990 77.340 ;
        RECT 71.690 76.490 71.990 77.340 ;
        RECT 73.690 76.490 73.990 77.340 ;
        RECT 87.125 76.490 87.425 77.340 ;
        RECT 89.125 76.490 89.425 77.340 ;
        RECT 91.125 76.490 91.425 77.340 ;
        RECT 93.125 76.490 93.425 77.340 ;
        RECT 95.125 76.490 95.425 77.340 ;
        RECT 97.125 76.490 97.425 77.340 ;
        RECT 99.125 76.490 99.425 77.340 ;
        RECT 101.125 76.490 101.425 77.340 ;
        RECT 103.125 76.490 103.425 77.340 ;
        RECT 105.125 76.490 105.425 77.340 ;
        RECT 107.125 76.490 107.425 77.340 ;
        RECT 109.125 76.490 109.425 77.340 ;
        RECT 111.125 76.490 111.425 77.340 ;
        RECT 113.125 76.490 113.425 77.340 ;
        RECT 115.125 76.490 115.425 77.340 ;
        RECT 117.125 76.490 117.425 77.340 ;
        RECT 119.125 76.490 119.425 77.340 ;
        RECT 121.125 76.490 121.425 77.340 ;
        RECT 123.125 76.490 123.425 77.340 ;
        RECT 125.125 76.490 125.425 77.340 ;
        RECT 127.125 76.490 127.425 77.340 ;
        RECT 129.125 76.490 129.425 77.340 ;
        RECT 131.125 76.490 131.425 77.340 ;
        RECT 133.125 76.490 133.425 77.340 ;
        RECT 135.125 76.490 135.425 77.340 ;
        RECT 137.125 76.490 137.425 77.340 ;
        RECT 139.125 76.490 139.425 77.340 ;
        RECT 141.125 76.490 141.425 77.340 ;
        RECT 143.125 76.490 143.425 77.340 ;
        RECT 145.125 76.490 145.425 77.340 ;
        RECT 147.125 76.490 147.425 77.340 ;
        RECT 149.125 76.490 149.425 77.340 ;
        RECT 151.125 76.490 151.425 77.340 ;
        RECT 153.125 76.490 153.425 77.340 ;
        RECT 7.340 75.490 8.340 76.490 ;
        RECT 9.340 75.490 10.340 76.490 ;
        RECT 11.340 75.490 12.340 76.490 ;
        RECT 13.340 75.490 14.340 76.490 ;
        RECT 15.340 75.490 16.340 76.490 ;
        RECT 17.340 75.490 18.340 76.490 ;
        RECT 19.340 75.490 20.340 76.490 ;
        RECT 21.340 75.490 22.340 76.490 ;
        RECT 23.340 75.490 24.340 76.490 ;
        RECT 25.340 75.490 26.340 76.490 ;
        RECT 27.340 75.490 28.340 76.490 ;
        RECT 29.340 75.490 30.340 76.490 ;
        RECT 31.340 75.490 32.340 76.490 ;
        RECT 33.340 75.490 34.340 76.490 ;
        RECT 35.340 75.490 36.340 76.490 ;
        RECT 37.340 75.490 38.340 76.490 ;
        RECT 39.340 75.490 40.340 76.490 ;
        RECT 41.340 75.490 42.340 76.490 ;
        RECT 43.340 75.490 44.340 76.490 ;
        RECT 45.340 75.490 46.340 76.490 ;
        RECT 47.340 75.490 48.340 76.490 ;
        RECT 49.340 75.490 50.340 76.490 ;
        RECT 51.340 75.490 52.340 76.490 ;
        RECT 53.340 75.490 54.340 76.490 ;
        RECT 55.340 75.490 56.340 76.490 ;
        RECT 57.340 75.490 58.340 76.490 ;
        RECT 59.340 75.490 60.340 76.490 ;
        RECT 61.340 75.490 62.340 76.490 ;
        RECT 63.340 75.490 64.340 76.490 ;
        RECT 65.340 75.490 66.340 76.490 ;
        RECT 67.340 75.490 68.340 76.490 ;
        RECT 69.340 75.490 70.340 76.490 ;
        RECT 71.340 75.490 72.340 76.490 ;
        RECT 73.340 75.490 74.340 76.490 ;
        RECT 86.775 75.490 87.775 76.490 ;
        RECT 88.775 75.490 89.775 76.490 ;
        RECT 90.775 75.490 91.775 76.490 ;
        RECT 92.775 75.490 93.775 76.490 ;
        RECT 94.775 75.490 95.775 76.490 ;
        RECT 96.775 75.490 97.775 76.490 ;
        RECT 98.775 75.490 99.775 76.490 ;
        RECT 100.775 75.490 101.775 76.490 ;
        RECT 102.775 75.490 103.775 76.490 ;
        RECT 104.775 75.490 105.775 76.490 ;
        RECT 106.775 75.490 107.775 76.490 ;
        RECT 108.775 75.490 109.775 76.490 ;
        RECT 110.775 75.490 111.775 76.490 ;
        RECT 112.775 75.490 113.775 76.490 ;
        RECT 114.775 75.490 115.775 76.490 ;
        RECT 116.775 75.490 117.775 76.490 ;
        RECT 118.775 75.490 119.775 76.490 ;
        RECT 120.775 75.490 121.775 76.490 ;
        RECT 122.775 75.490 123.775 76.490 ;
        RECT 124.775 75.490 125.775 76.490 ;
        RECT 126.775 75.490 127.775 76.490 ;
        RECT 128.775 75.490 129.775 76.490 ;
        RECT 130.775 75.490 131.775 76.490 ;
        RECT 132.775 75.490 133.775 76.490 ;
        RECT 134.775 75.490 135.775 76.490 ;
        RECT 136.775 75.490 137.775 76.490 ;
        RECT 138.775 75.490 139.775 76.490 ;
        RECT 140.775 75.490 141.775 76.490 ;
        RECT 142.775 75.490 143.775 76.490 ;
        RECT 144.775 75.490 145.775 76.490 ;
        RECT 146.775 75.490 147.775 76.490 ;
        RECT 148.775 75.490 149.775 76.490 ;
        RECT 150.775 75.490 151.775 76.490 ;
        RECT 152.775 75.490 153.775 76.490 ;
        RECT 7.690 74.640 7.990 75.490 ;
        RECT 9.690 74.640 9.990 75.490 ;
        RECT 11.690 74.640 11.990 75.490 ;
        RECT 13.690 74.640 13.990 75.490 ;
        RECT 15.690 74.640 15.990 75.490 ;
        RECT 17.690 74.640 17.990 75.490 ;
        RECT 19.690 74.640 19.990 75.490 ;
        RECT 21.690 74.640 21.990 75.490 ;
        RECT 23.690 74.640 23.990 75.490 ;
        RECT 25.690 74.640 25.990 75.490 ;
        RECT 27.690 74.640 27.990 75.490 ;
        RECT 29.690 74.640 29.990 75.490 ;
        RECT 31.690 74.640 31.990 75.490 ;
        RECT 33.690 74.640 33.990 75.490 ;
        RECT 35.690 74.640 35.990 75.490 ;
        RECT 37.690 74.640 37.990 75.490 ;
        RECT 39.690 74.640 39.990 75.490 ;
        RECT 41.690 74.640 41.990 75.490 ;
        RECT 43.690 74.640 43.990 75.490 ;
        RECT 45.690 74.640 45.990 75.490 ;
        RECT 47.690 74.640 47.990 75.490 ;
        RECT 49.690 74.640 49.990 75.490 ;
        RECT 51.690 74.640 51.990 75.490 ;
        RECT 53.690 74.640 53.990 75.490 ;
        RECT 55.690 74.640 55.990 75.490 ;
        RECT 57.690 74.640 57.990 75.490 ;
        RECT 59.690 74.640 59.990 75.490 ;
        RECT 61.690 74.640 61.990 75.490 ;
        RECT 63.690 74.640 63.990 75.490 ;
        RECT 65.690 74.640 65.990 75.490 ;
        RECT 67.690 74.640 67.990 75.490 ;
        RECT 69.690 74.640 69.990 75.490 ;
        RECT 71.690 74.640 71.990 75.490 ;
        RECT 73.690 74.640 73.990 75.490 ;
        RECT 87.125 74.640 87.425 75.490 ;
        RECT 89.125 74.640 89.425 75.490 ;
        RECT 91.125 74.640 91.425 75.490 ;
        RECT 93.125 74.640 93.425 75.490 ;
        RECT 95.125 74.640 95.425 75.490 ;
        RECT 97.125 74.640 97.425 75.490 ;
        RECT 99.125 74.640 99.425 75.490 ;
        RECT 101.125 74.640 101.425 75.490 ;
        RECT 103.125 74.640 103.425 75.490 ;
        RECT 105.125 74.640 105.425 75.490 ;
        RECT 107.125 74.640 107.425 75.490 ;
        RECT 109.125 74.640 109.425 75.490 ;
        RECT 111.125 74.640 111.425 75.490 ;
        RECT 113.125 74.640 113.425 75.490 ;
        RECT 115.125 74.640 115.425 75.490 ;
        RECT 117.125 74.640 117.425 75.490 ;
        RECT 119.125 74.640 119.425 75.490 ;
        RECT 121.125 74.640 121.425 75.490 ;
        RECT 123.125 74.640 123.425 75.490 ;
        RECT 125.125 74.640 125.425 75.490 ;
        RECT 127.125 74.640 127.425 75.490 ;
        RECT 129.125 74.640 129.425 75.490 ;
        RECT 131.125 74.640 131.425 75.490 ;
        RECT 133.125 74.640 133.425 75.490 ;
        RECT 135.125 74.640 135.425 75.490 ;
        RECT 137.125 74.640 137.425 75.490 ;
        RECT 139.125 74.640 139.425 75.490 ;
        RECT 141.125 74.640 141.425 75.490 ;
        RECT 143.125 74.640 143.425 75.490 ;
        RECT 145.125 74.640 145.425 75.490 ;
        RECT 147.125 74.640 147.425 75.490 ;
        RECT 149.125 74.640 149.425 75.490 ;
        RECT 151.125 74.640 151.425 75.490 ;
        RECT 153.125 74.640 153.425 75.490 ;
        RECT 7.340 73.640 8.340 74.640 ;
        RECT 9.340 73.640 10.340 74.640 ;
        RECT 11.340 73.640 12.340 74.640 ;
        RECT 13.340 73.640 14.340 74.640 ;
        RECT 15.340 73.640 16.340 74.640 ;
        RECT 17.340 73.640 18.340 74.640 ;
        RECT 19.340 73.640 20.340 74.640 ;
        RECT 21.340 73.640 22.340 74.640 ;
        RECT 23.340 73.640 24.340 74.640 ;
        RECT 25.340 73.640 26.340 74.640 ;
        RECT 27.340 73.640 28.340 74.640 ;
        RECT 29.340 73.640 30.340 74.640 ;
        RECT 31.340 73.640 32.340 74.640 ;
        RECT 33.340 73.640 34.340 74.640 ;
        RECT 35.340 73.640 36.340 74.640 ;
        RECT 37.340 73.640 38.340 74.640 ;
        RECT 39.340 73.640 40.340 74.640 ;
        RECT 41.340 73.640 42.340 74.640 ;
        RECT 43.340 73.640 44.340 74.640 ;
        RECT 45.340 73.640 46.340 74.640 ;
        RECT 47.340 73.640 48.340 74.640 ;
        RECT 49.340 73.640 50.340 74.640 ;
        RECT 51.340 73.640 52.340 74.640 ;
        RECT 53.340 73.640 54.340 74.640 ;
        RECT 55.340 73.640 56.340 74.640 ;
        RECT 57.340 73.640 58.340 74.640 ;
        RECT 59.340 73.640 60.340 74.640 ;
        RECT 61.340 73.640 62.340 74.640 ;
        RECT 63.340 73.640 64.340 74.640 ;
        RECT 65.340 73.640 66.340 74.640 ;
        RECT 67.340 73.640 68.340 74.640 ;
        RECT 69.340 73.640 70.340 74.640 ;
        RECT 71.340 73.640 72.340 74.640 ;
        RECT 73.340 73.640 74.340 74.640 ;
        RECT 86.775 73.640 87.775 74.640 ;
        RECT 88.775 73.640 89.775 74.640 ;
        RECT 90.775 73.640 91.775 74.640 ;
        RECT 92.775 73.640 93.775 74.640 ;
        RECT 94.775 73.640 95.775 74.640 ;
        RECT 96.775 73.640 97.775 74.640 ;
        RECT 98.775 73.640 99.775 74.640 ;
        RECT 100.775 73.640 101.775 74.640 ;
        RECT 102.775 73.640 103.775 74.640 ;
        RECT 104.775 73.640 105.775 74.640 ;
        RECT 106.775 73.640 107.775 74.640 ;
        RECT 108.775 73.640 109.775 74.640 ;
        RECT 110.775 73.640 111.775 74.640 ;
        RECT 112.775 73.640 113.775 74.640 ;
        RECT 114.775 73.640 115.775 74.640 ;
        RECT 116.775 73.640 117.775 74.640 ;
        RECT 118.775 73.640 119.775 74.640 ;
        RECT 120.775 73.640 121.775 74.640 ;
        RECT 122.775 73.640 123.775 74.640 ;
        RECT 124.775 73.640 125.775 74.640 ;
        RECT 126.775 73.640 127.775 74.640 ;
        RECT 128.775 73.640 129.775 74.640 ;
        RECT 130.775 73.640 131.775 74.640 ;
        RECT 132.775 73.640 133.775 74.640 ;
        RECT 134.775 73.640 135.775 74.640 ;
        RECT 136.775 73.640 137.775 74.640 ;
        RECT 138.775 73.640 139.775 74.640 ;
        RECT 140.775 73.640 141.775 74.640 ;
        RECT 142.775 73.640 143.775 74.640 ;
        RECT 144.775 73.640 145.775 74.640 ;
        RECT 146.775 73.640 147.775 74.640 ;
        RECT 148.775 73.640 149.775 74.640 ;
        RECT 150.775 73.640 151.775 74.640 ;
        RECT 152.775 73.640 153.775 74.640 ;
        RECT 7.690 72.790 7.990 73.640 ;
        RECT 9.690 72.790 9.990 73.640 ;
        RECT 11.690 72.790 11.990 73.640 ;
        RECT 13.690 72.790 13.990 73.640 ;
        RECT 15.690 72.790 15.990 73.640 ;
        RECT 17.690 72.790 17.990 73.640 ;
        RECT 19.690 72.790 19.990 73.640 ;
        RECT 21.690 72.790 21.990 73.640 ;
        RECT 23.690 72.790 23.990 73.640 ;
        RECT 25.690 72.790 25.990 73.640 ;
        RECT 27.690 72.790 27.990 73.640 ;
        RECT 29.690 72.790 29.990 73.640 ;
        RECT 31.690 72.790 31.990 73.640 ;
        RECT 33.690 72.790 33.990 73.640 ;
        RECT 35.690 72.790 35.990 73.640 ;
        RECT 37.690 72.790 37.990 73.640 ;
        RECT 39.690 72.790 39.990 73.640 ;
        RECT 41.690 72.790 41.990 73.640 ;
        RECT 43.690 72.790 43.990 73.640 ;
        RECT 45.690 72.790 45.990 73.640 ;
        RECT 47.690 72.790 47.990 73.640 ;
        RECT 49.690 72.790 49.990 73.640 ;
        RECT 51.690 72.790 51.990 73.640 ;
        RECT 53.690 72.790 53.990 73.640 ;
        RECT 55.690 72.790 55.990 73.640 ;
        RECT 57.690 72.790 57.990 73.640 ;
        RECT 59.690 72.790 59.990 73.640 ;
        RECT 61.690 72.790 61.990 73.640 ;
        RECT 63.690 72.790 63.990 73.640 ;
        RECT 65.690 72.790 65.990 73.640 ;
        RECT 67.690 72.790 67.990 73.640 ;
        RECT 69.690 72.790 69.990 73.640 ;
        RECT 71.690 72.790 71.990 73.640 ;
        RECT 73.690 72.790 73.990 73.640 ;
        RECT 87.125 72.790 87.425 73.640 ;
        RECT 89.125 72.790 89.425 73.640 ;
        RECT 91.125 72.790 91.425 73.640 ;
        RECT 93.125 72.790 93.425 73.640 ;
        RECT 95.125 72.790 95.425 73.640 ;
        RECT 97.125 72.790 97.425 73.640 ;
        RECT 99.125 72.790 99.425 73.640 ;
        RECT 101.125 72.790 101.425 73.640 ;
        RECT 103.125 72.790 103.425 73.640 ;
        RECT 105.125 72.790 105.425 73.640 ;
        RECT 107.125 72.790 107.425 73.640 ;
        RECT 109.125 72.790 109.425 73.640 ;
        RECT 111.125 72.790 111.425 73.640 ;
        RECT 113.125 72.790 113.425 73.640 ;
        RECT 115.125 72.790 115.425 73.640 ;
        RECT 117.125 72.790 117.425 73.640 ;
        RECT 119.125 72.790 119.425 73.640 ;
        RECT 121.125 72.790 121.425 73.640 ;
        RECT 123.125 72.790 123.425 73.640 ;
        RECT 125.125 72.790 125.425 73.640 ;
        RECT 127.125 72.790 127.425 73.640 ;
        RECT 129.125 72.790 129.425 73.640 ;
        RECT 131.125 72.790 131.425 73.640 ;
        RECT 133.125 72.790 133.425 73.640 ;
        RECT 135.125 72.790 135.425 73.640 ;
        RECT 137.125 72.790 137.425 73.640 ;
        RECT 139.125 72.790 139.425 73.640 ;
        RECT 141.125 72.790 141.425 73.640 ;
        RECT 143.125 72.790 143.425 73.640 ;
        RECT 145.125 72.790 145.425 73.640 ;
        RECT 147.125 72.790 147.425 73.640 ;
        RECT 149.125 72.790 149.425 73.640 ;
        RECT 151.125 72.790 151.425 73.640 ;
        RECT 153.125 72.790 153.425 73.640 ;
        RECT 7.340 71.790 8.340 72.790 ;
        RECT 9.340 71.790 10.340 72.790 ;
        RECT 11.340 71.790 12.340 72.790 ;
        RECT 13.340 71.790 14.340 72.790 ;
        RECT 15.340 71.790 16.340 72.790 ;
        RECT 17.340 71.790 18.340 72.790 ;
        RECT 19.340 71.790 20.340 72.790 ;
        RECT 21.340 71.790 22.340 72.790 ;
        RECT 23.340 71.790 24.340 72.790 ;
        RECT 25.340 71.790 26.340 72.790 ;
        RECT 27.340 71.790 28.340 72.790 ;
        RECT 29.340 71.790 30.340 72.790 ;
        RECT 31.340 71.790 32.340 72.790 ;
        RECT 33.340 71.790 34.340 72.790 ;
        RECT 35.340 71.790 36.340 72.790 ;
        RECT 37.340 71.790 38.340 72.790 ;
        RECT 39.340 71.790 40.340 72.790 ;
        RECT 41.340 71.790 42.340 72.790 ;
        RECT 43.340 71.790 44.340 72.790 ;
        RECT 45.340 71.790 46.340 72.790 ;
        RECT 47.340 71.790 48.340 72.790 ;
        RECT 49.340 71.790 50.340 72.790 ;
        RECT 51.340 71.790 52.340 72.790 ;
        RECT 53.340 71.790 54.340 72.790 ;
        RECT 55.340 71.790 56.340 72.790 ;
        RECT 57.340 71.790 58.340 72.790 ;
        RECT 59.340 71.790 60.340 72.790 ;
        RECT 61.340 71.790 62.340 72.790 ;
        RECT 63.340 71.790 64.340 72.790 ;
        RECT 65.340 71.790 66.340 72.790 ;
        RECT 67.340 71.790 68.340 72.790 ;
        RECT 69.340 71.790 70.340 72.790 ;
        RECT 71.340 71.790 72.340 72.790 ;
        RECT 73.340 71.790 74.340 72.790 ;
        RECT 86.775 71.790 87.775 72.790 ;
        RECT 88.775 71.790 89.775 72.790 ;
        RECT 90.775 71.790 91.775 72.790 ;
        RECT 92.775 71.790 93.775 72.790 ;
        RECT 94.775 71.790 95.775 72.790 ;
        RECT 96.775 71.790 97.775 72.790 ;
        RECT 98.775 71.790 99.775 72.790 ;
        RECT 100.775 71.790 101.775 72.790 ;
        RECT 102.775 71.790 103.775 72.790 ;
        RECT 104.775 71.790 105.775 72.790 ;
        RECT 106.775 71.790 107.775 72.790 ;
        RECT 108.775 71.790 109.775 72.790 ;
        RECT 110.775 71.790 111.775 72.790 ;
        RECT 112.775 71.790 113.775 72.790 ;
        RECT 114.775 71.790 115.775 72.790 ;
        RECT 116.775 71.790 117.775 72.790 ;
        RECT 118.775 71.790 119.775 72.790 ;
        RECT 120.775 71.790 121.775 72.790 ;
        RECT 122.775 71.790 123.775 72.790 ;
        RECT 124.775 71.790 125.775 72.790 ;
        RECT 126.775 71.790 127.775 72.790 ;
        RECT 128.775 71.790 129.775 72.790 ;
        RECT 130.775 71.790 131.775 72.790 ;
        RECT 132.775 71.790 133.775 72.790 ;
        RECT 134.775 71.790 135.775 72.790 ;
        RECT 136.775 71.790 137.775 72.790 ;
        RECT 138.775 71.790 139.775 72.790 ;
        RECT 140.775 71.790 141.775 72.790 ;
        RECT 142.775 71.790 143.775 72.790 ;
        RECT 144.775 71.790 145.775 72.790 ;
        RECT 146.775 71.790 147.775 72.790 ;
        RECT 148.775 71.790 149.775 72.790 ;
        RECT 150.775 71.790 151.775 72.790 ;
        RECT 152.775 71.790 153.775 72.790 ;
        RECT 7.690 70.940 7.990 71.790 ;
        RECT 9.690 70.940 9.990 71.790 ;
        RECT 11.690 70.940 11.990 71.790 ;
        RECT 13.690 70.940 13.990 71.790 ;
        RECT 15.690 70.940 15.990 71.790 ;
        RECT 17.690 70.940 17.990 71.790 ;
        RECT 19.690 70.940 19.990 71.790 ;
        RECT 21.690 70.940 21.990 71.790 ;
        RECT 23.690 70.940 23.990 71.790 ;
        RECT 25.690 70.940 25.990 71.790 ;
        RECT 27.690 70.940 27.990 71.790 ;
        RECT 29.690 70.940 29.990 71.790 ;
        RECT 31.690 70.940 31.990 71.790 ;
        RECT 33.690 70.940 33.990 71.790 ;
        RECT 35.690 70.940 35.990 71.790 ;
        RECT 37.690 70.940 37.990 71.790 ;
        RECT 39.690 70.940 39.990 71.790 ;
        RECT 41.690 70.940 41.990 71.790 ;
        RECT 43.690 70.940 43.990 71.790 ;
        RECT 45.690 70.940 45.990 71.790 ;
        RECT 47.690 70.940 47.990 71.790 ;
        RECT 49.690 70.940 49.990 71.790 ;
        RECT 51.690 70.940 51.990 71.790 ;
        RECT 53.690 70.940 53.990 71.790 ;
        RECT 55.690 70.940 55.990 71.790 ;
        RECT 57.690 70.940 57.990 71.790 ;
        RECT 59.690 70.940 59.990 71.790 ;
        RECT 61.690 70.940 61.990 71.790 ;
        RECT 63.690 70.940 63.990 71.790 ;
        RECT 65.690 70.940 65.990 71.790 ;
        RECT 67.690 70.940 67.990 71.790 ;
        RECT 69.690 70.940 69.990 71.790 ;
        RECT 71.690 70.940 71.990 71.790 ;
        RECT 73.690 70.940 73.990 71.790 ;
        RECT 87.125 70.940 87.425 71.790 ;
        RECT 89.125 70.940 89.425 71.790 ;
        RECT 91.125 70.940 91.425 71.790 ;
        RECT 93.125 70.940 93.425 71.790 ;
        RECT 95.125 70.940 95.425 71.790 ;
        RECT 97.125 70.940 97.425 71.790 ;
        RECT 99.125 70.940 99.425 71.790 ;
        RECT 101.125 70.940 101.425 71.790 ;
        RECT 103.125 70.940 103.425 71.790 ;
        RECT 105.125 70.940 105.425 71.790 ;
        RECT 107.125 70.940 107.425 71.790 ;
        RECT 109.125 70.940 109.425 71.790 ;
        RECT 111.125 70.940 111.425 71.790 ;
        RECT 113.125 70.940 113.425 71.790 ;
        RECT 115.125 70.940 115.425 71.790 ;
        RECT 117.125 70.940 117.425 71.790 ;
        RECT 119.125 70.940 119.425 71.790 ;
        RECT 121.125 70.940 121.425 71.790 ;
        RECT 123.125 70.940 123.425 71.790 ;
        RECT 125.125 70.940 125.425 71.790 ;
        RECT 127.125 70.940 127.425 71.790 ;
        RECT 129.125 70.940 129.425 71.790 ;
        RECT 131.125 70.940 131.425 71.790 ;
        RECT 133.125 70.940 133.425 71.790 ;
        RECT 135.125 70.940 135.425 71.790 ;
        RECT 137.125 70.940 137.425 71.790 ;
        RECT 139.125 70.940 139.425 71.790 ;
        RECT 141.125 70.940 141.425 71.790 ;
        RECT 143.125 70.940 143.425 71.790 ;
        RECT 145.125 70.940 145.425 71.790 ;
        RECT 147.125 70.940 147.425 71.790 ;
        RECT 149.125 70.940 149.425 71.790 ;
        RECT 151.125 70.940 151.425 71.790 ;
        RECT 153.125 70.940 153.425 71.790 ;
        RECT 7.340 69.940 8.340 70.940 ;
        RECT 9.340 69.940 10.340 70.940 ;
        RECT 11.340 69.940 12.340 70.940 ;
        RECT 13.340 69.940 14.340 70.940 ;
        RECT 15.340 69.940 16.340 70.940 ;
        RECT 17.340 69.940 18.340 70.940 ;
        RECT 19.340 69.940 20.340 70.940 ;
        RECT 21.340 69.940 22.340 70.940 ;
        RECT 23.340 69.940 24.340 70.940 ;
        RECT 25.340 69.940 26.340 70.940 ;
        RECT 27.340 69.940 28.340 70.940 ;
        RECT 29.340 69.940 30.340 70.940 ;
        RECT 31.340 69.940 32.340 70.940 ;
        RECT 33.340 69.940 34.340 70.940 ;
        RECT 35.340 69.940 36.340 70.940 ;
        RECT 37.340 69.940 38.340 70.940 ;
        RECT 39.340 69.940 40.340 70.940 ;
        RECT 41.340 69.940 42.340 70.940 ;
        RECT 43.340 69.940 44.340 70.940 ;
        RECT 45.340 69.940 46.340 70.940 ;
        RECT 47.340 69.940 48.340 70.940 ;
        RECT 49.340 69.940 50.340 70.940 ;
        RECT 51.340 69.940 52.340 70.940 ;
        RECT 53.340 69.940 54.340 70.940 ;
        RECT 55.340 69.940 56.340 70.940 ;
        RECT 57.340 69.940 58.340 70.940 ;
        RECT 59.340 69.940 60.340 70.940 ;
        RECT 61.340 69.940 62.340 70.940 ;
        RECT 63.340 69.940 64.340 70.940 ;
        RECT 65.340 69.940 66.340 70.940 ;
        RECT 67.340 69.940 68.340 70.940 ;
        RECT 69.340 69.940 70.340 70.940 ;
        RECT 71.340 69.940 72.340 70.940 ;
        RECT 73.340 69.940 74.340 70.940 ;
        RECT 86.775 69.940 87.775 70.940 ;
        RECT 88.775 69.940 89.775 70.940 ;
        RECT 90.775 69.940 91.775 70.940 ;
        RECT 92.775 69.940 93.775 70.940 ;
        RECT 94.775 69.940 95.775 70.940 ;
        RECT 96.775 69.940 97.775 70.940 ;
        RECT 98.775 69.940 99.775 70.940 ;
        RECT 100.775 69.940 101.775 70.940 ;
        RECT 102.775 69.940 103.775 70.940 ;
        RECT 104.775 69.940 105.775 70.940 ;
        RECT 106.775 69.940 107.775 70.940 ;
        RECT 108.775 69.940 109.775 70.940 ;
        RECT 110.775 69.940 111.775 70.940 ;
        RECT 112.775 69.940 113.775 70.940 ;
        RECT 114.775 69.940 115.775 70.940 ;
        RECT 116.775 69.940 117.775 70.940 ;
        RECT 118.775 69.940 119.775 70.940 ;
        RECT 120.775 69.940 121.775 70.940 ;
        RECT 122.775 69.940 123.775 70.940 ;
        RECT 124.775 69.940 125.775 70.940 ;
        RECT 126.775 69.940 127.775 70.940 ;
        RECT 128.775 69.940 129.775 70.940 ;
        RECT 130.775 69.940 131.775 70.940 ;
        RECT 132.775 69.940 133.775 70.940 ;
        RECT 134.775 69.940 135.775 70.940 ;
        RECT 136.775 69.940 137.775 70.940 ;
        RECT 138.775 69.940 139.775 70.940 ;
        RECT 140.775 69.940 141.775 70.940 ;
        RECT 142.775 69.940 143.775 70.940 ;
        RECT 144.775 69.940 145.775 70.940 ;
        RECT 146.775 69.940 147.775 70.940 ;
        RECT 148.775 69.940 149.775 70.940 ;
        RECT 150.775 69.940 151.775 70.940 ;
        RECT 152.775 69.940 153.775 70.940 ;
        RECT 7.690 69.090 7.990 69.940 ;
        RECT 9.690 69.090 9.990 69.940 ;
        RECT 11.690 69.090 11.990 69.940 ;
        RECT 13.690 69.090 13.990 69.940 ;
        RECT 15.690 69.090 15.990 69.940 ;
        RECT 17.690 69.090 17.990 69.940 ;
        RECT 19.690 69.090 19.990 69.940 ;
        RECT 21.690 69.090 21.990 69.940 ;
        RECT 23.690 69.090 23.990 69.940 ;
        RECT 25.690 69.090 25.990 69.940 ;
        RECT 27.690 69.090 27.990 69.940 ;
        RECT 29.690 69.090 29.990 69.940 ;
        RECT 31.690 69.090 31.990 69.940 ;
        RECT 33.690 69.090 33.990 69.940 ;
        RECT 35.690 69.090 35.990 69.940 ;
        RECT 37.690 69.090 37.990 69.940 ;
        RECT 39.690 69.090 39.990 69.940 ;
        RECT 41.690 69.090 41.990 69.940 ;
        RECT 43.690 69.090 43.990 69.940 ;
        RECT 45.690 69.090 45.990 69.940 ;
        RECT 47.690 69.090 47.990 69.940 ;
        RECT 49.690 69.090 49.990 69.940 ;
        RECT 51.690 69.090 51.990 69.940 ;
        RECT 53.690 69.090 53.990 69.940 ;
        RECT 55.690 69.090 55.990 69.940 ;
        RECT 57.690 69.090 57.990 69.940 ;
        RECT 59.690 69.090 59.990 69.940 ;
        RECT 61.690 69.090 61.990 69.940 ;
        RECT 63.690 69.090 63.990 69.940 ;
        RECT 65.690 69.090 65.990 69.940 ;
        RECT 67.690 69.090 67.990 69.940 ;
        RECT 69.690 69.090 69.990 69.940 ;
        RECT 71.690 69.090 71.990 69.940 ;
        RECT 73.690 69.090 73.990 69.940 ;
        RECT 87.125 69.090 87.425 69.940 ;
        RECT 89.125 69.090 89.425 69.940 ;
        RECT 91.125 69.090 91.425 69.940 ;
        RECT 93.125 69.090 93.425 69.940 ;
        RECT 95.125 69.090 95.425 69.940 ;
        RECT 97.125 69.090 97.425 69.940 ;
        RECT 99.125 69.090 99.425 69.940 ;
        RECT 101.125 69.090 101.425 69.940 ;
        RECT 103.125 69.090 103.425 69.940 ;
        RECT 105.125 69.090 105.425 69.940 ;
        RECT 107.125 69.090 107.425 69.940 ;
        RECT 109.125 69.090 109.425 69.940 ;
        RECT 111.125 69.090 111.425 69.940 ;
        RECT 113.125 69.090 113.425 69.940 ;
        RECT 115.125 69.090 115.425 69.940 ;
        RECT 117.125 69.090 117.425 69.940 ;
        RECT 119.125 69.090 119.425 69.940 ;
        RECT 121.125 69.090 121.425 69.940 ;
        RECT 123.125 69.090 123.425 69.940 ;
        RECT 125.125 69.090 125.425 69.940 ;
        RECT 127.125 69.090 127.425 69.940 ;
        RECT 129.125 69.090 129.425 69.940 ;
        RECT 131.125 69.090 131.425 69.940 ;
        RECT 133.125 69.090 133.425 69.940 ;
        RECT 135.125 69.090 135.425 69.940 ;
        RECT 137.125 69.090 137.425 69.940 ;
        RECT 139.125 69.090 139.425 69.940 ;
        RECT 141.125 69.090 141.425 69.940 ;
        RECT 143.125 69.090 143.425 69.940 ;
        RECT 145.125 69.090 145.425 69.940 ;
        RECT 147.125 69.090 147.425 69.940 ;
        RECT 149.125 69.090 149.425 69.940 ;
        RECT 151.125 69.090 151.425 69.940 ;
        RECT 153.125 69.090 153.425 69.940 ;
        RECT 7.340 68.090 8.340 69.090 ;
        RECT 9.340 68.090 10.340 69.090 ;
        RECT 11.340 68.090 12.340 69.090 ;
        RECT 13.340 68.090 14.340 69.090 ;
        RECT 15.340 68.090 16.340 69.090 ;
        RECT 17.340 68.090 18.340 69.090 ;
        RECT 19.340 68.090 20.340 69.090 ;
        RECT 21.340 68.090 22.340 69.090 ;
        RECT 23.340 68.090 24.340 69.090 ;
        RECT 25.340 68.090 26.340 69.090 ;
        RECT 27.340 68.090 28.340 69.090 ;
        RECT 29.340 68.090 30.340 69.090 ;
        RECT 31.340 68.090 32.340 69.090 ;
        RECT 33.340 68.090 34.340 69.090 ;
        RECT 35.340 68.090 36.340 69.090 ;
        RECT 37.340 68.090 38.340 69.090 ;
        RECT 39.340 68.090 40.340 69.090 ;
        RECT 41.340 68.090 42.340 69.090 ;
        RECT 43.340 68.090 44.340 69.090 ;
        RECT 45.340 68.090 46.340 69.090 ;
        RECT 47.340 68.090 48.340 69.090 ;
        RECT 49.340 68.090 50.340 69.090 ;
        RECT 51.340 68.090 52.340 69.090 ;
        RECT 53.340 68.090 54.340 69.090 ;
        RECT 55.340 68.090 56.340 69.090 ;
        RECT 57.340 68.090 58.340 69.090 ;
        RECT 59.340 68.090 60.340 69.090 ;
        RECT 61.340 68.090 62.340 69.090 ;
        RECT 63.340 68.090 64.340 69.090 ;
        RECT 65.340 68.090 66.340 69.090 ;
        RECT 67.340 68.090 68.340 69.090 ;
        RECT 69.340 68.090 70.340 69.090 ;
        RECT 71.340 68.090 72.340 69.090 ;
        RECT 73.340 68.090 74.340 69.090 ;
        RECT 86.775 68.090 87.775 69.090 ;
        RECT 88.775 68.090 89.775 69.090 ;
        RECT 90.775 68.090 91.775 69.090 ;
        RECT 92.775 68.090 93.775 69.090 ;
        RECT 94.775 68.090 95.775 69.090 ;
        RECT 96.775 68.090 97.775 69.090 ;
        RECT 98.775 68.090 99.775 69.090 ;
        RECT 100.775 68.090 101.775 69.090 ;
        RECT 102.775 68.090 103.775 69.090 ;
        RECT 104.775 68.090 105.775 69.090 ;
        RECT 106.775 68.090 107.775 69.090 ;
        RECT 108.775 68.090 109.775 69.090 ;
        RECT 110.775 68.090 111.775 69.090 ;
        RECT 112.775 68.090 113.775 69.090 ;
        RECT 114.775 68.090 115.775 69.090 ;
        RECT 116.775 68.090 117.775 69.090 ;
        RECT 118.775 68.090 119.775 69.090 ;
        RECT 120.775 68.090 121.775 69.090 ;
        RECT 122.775 68.090 123.775 69.090 ;
        RECT 124.775 68.090 125.775 69.090 ;
        RECT 126.775 68.090 127.775 69.090 ;
        RECT 128.775 68.090 129.775 69.090 ;
        RECT 130.775 68.090 131.775 69.090 ;
        RECT 132.775 68.090 133.775 69.090 ;
        RECT 134.775 68.090 135.775 69.090 ;
        RECT 136.775 68.090 137.775 69.090 ;
        RECT 138.775 68.090 139.775 69.090 ;
        RECT 140.775 68.090 141.775 69.090 ;
        RECT 142.775 68.090 143.775 69.090 ;
        RECT 144.775 68.090 145.775 69.090 ;
        RECT 146.775 68.090 147.775 69.090 ;
        RECT 148.775 68.090 149.775 69.090 ;
        RECT 150.775 68.090 151.775 69.090 ;
        RECT 152.775 68.090 153.775 69.090 ;
        RECT 7.690 67.240 7.990 68.090 ;
        RECT 9.690 67.240 9.990 68.090 ;
        RECT 11.690 67.240 11.990 68.090 ;
        RECT 13.690 67.240 13.990 68.090 ;
        RECT 15.690 67.240 15.990 68.090 ;
        RECT 17.690 67.240 17.990 68.090 ;
        RECT 19.690 67.240 19.990 68.090 ;
        RECT 21.690 67.240 21.990 68.090 ;
        RECT 23.690 67.240 23.990 68.090 ;
        RECT 25.690 67.240 25.990 68.090 ;
        RECT 27.690 67.240 27.990 68.090 ;
        RECT 29.690 67.240 29.990 68.090 ;
        RECT 31.690 67.240 31.990 68.090 ;
        RECT 33.690 67.240 33.990 68.090 ;
        RECT 35.690 67.240 35.990 68.090 ;
        RECT 37.690 67.240 37.990 68.090 ;
        RECT 39.690 67.240 39.990 68.090 ;
        RECT 41.690 67.240 41.990 68.090 ;
        RECT 43.690 67.240 43.990 68.090 ;
        RECT 45.690 67.240 45.990 68.090 ;
        RECT 47.690 67.240 47.990 68.090 ;
        RECT 49.690 67.240 49.990 68.090 ;
        RECT 51.690 67.240 51.990 68.090 ;
        RECT 53.690 67.240 53.990 68.090 ;
        RECT 55.690 67.240 55.990 68.090 ;
        RECT 57.690 67.240 57.990 68.090 ;
        RECT 59.690 67.240 59.990 68.090 ;
        RECT 61.690 67.240 61.990 68.090 ;
        RECT 63.690 67.240 63.990 68.090 ;
        RECT 65.690 67.240 65.990 68.090 ;
        RECT 67.690 67.240 67.990 68.090 ;
        RECT 69.690 67.240 69.990 68.090 ;
        RECT 71.690 67.240 71.990 68.090 ;
        RECT 73.690 67.240 73.990 68.090 ;
        RECT 87.125 67.240 87.425 68.090 ;
        RECT 89.125 67.240 89.425 68.090 ;
        RECT 91.125 67.240 91.425 68.090 ;
        RECT 93.125 67.240 93.425 68.090 ;
        RECT 95.125 67.240 95.425 68.090 ;
        RECT 97.125 67.240 97.425 68.090 ;
        RECT 99.125 67.240 99.425 68.090 ;
        RECT 101.125 67.240 101.425 68.090 ;
        RECT 103.125 67.240 103.425 68.090 ;
        RECT 105.125 67.240 105.425 68.090 ;
        RECT 107.125 67.240 107.425 68.090 ;
        RECT 109.125 67.240 109.425 68.090 ;
        RECT 111.125 67.240 111.425 68.090 ;
        RECT 113.125 67.240 113.425 68.090 ;
        RECT 115.125 67.240 115.425 68.090 ;
        RECT 117.125 67.240 117.425 68.090 ;
        RECT 119.125 67.240 119.425 68.090 ;
        RECT 121.125 67.240 121.425 68.090 ;
        RECT 123.125 67.240 123.425 68.090 ;
        RECT 125.125 67.240 125.425 68.090 ;
        RECT 127.125 67.240 127.425 68.090 ;
        RECT 129.125 67.240 129.425 68.090 ;
        RECT 131.125 67.240 131.425 68.090 ;
        RECT 133.125 67.240 133.425 68.090 ;
        RECT 135.125 67.240 135.425 68.090 ;
        RECT 137.125 67.240 137.425 68.090 ;
        RECT 139.125 67.240 139.425 68.090 ;
        RECT 141.125 67.240 141.425 68.090 ;
        RECT 143.125 67.240 143.425 68.090 ;
        RECT 145.125 67.240 145.425 68.090 ;
        RECT 147.125 67.240 147.425 68.090 ;
        RECT 149.125 67.240 149.425 68.090 ;
        RECT 151.125 67.240 151.425 68.090 ;
        RECT 153.125 67.240 153.425 68.090 ;
        RECT 7.340 66.240 8.340 67.240 ;
        RECT 9.340 66.240 10.340 67.240 ;
        RECT 11.340 66.240 12.340 67.240 ;
        RECT 13.340 66.240 14.340 67.240 ;
        RECT 15.340 66.240 16.340 67.240 ;
        RECT 17.340 66.240 18.340 67.240 ;
        RECT 19.340 66.240 20.340 67.240 ;
        RECT 21.340 66.240 22.340 67.240 ;
        RECT 23.340 66.240 24.340 67.240 ;
        RECT 25.340 66.240 26.340 67.240 ;
        RECT 27.340 66.240 28.340 67.240 ;
        RECT 29.340 66.240 30.340 67.240 ;
        RECT 31.340 66.240 32.340 67.240 ;
        RECT 33.340 66.240 34.340 67.240 ;
        RECT 35.340 66.240 36.340 67.240 ;
        RECT 37.340 66.240 38.340 67.240 ;
        RECT 39.340 66.240 40.340 67.240 ;
        RECT 41.340 66.240 42.340 67.240 ;
        RECT 43.340 66.240 44.340 67.240 ;
        RECT 45.340 66.240 46.340 67.240 ;
        RECT 47.340 66.240 48.340 67.240 ;
        RECT 49.340 66.240 50.340 67.240 ;
        RECT 51.340 66.240 52.340 67.240 ;
        RECT 53.340 66.240 54.340 67.240 ;
        RECT 55.340 66.240 56.340 67.240 ;
        RECT 57.340 66.240 58.340 67.240 ;
        RECT 59.340 66.240 60.340 67.240 ;
        RECT 61.340 66.240 62.340 67.240 ;
        RECT 63.340 66.240 64.340 67.240 ;
        RECT 65.340 66.240 66.340 67.240 ;
        RECT 67.340 66.240 68.340 67.240 ;
        RECT 69.340 66.240 70.340 67.240 ;
        RECT 71.340 66.240 72.340 67.240 ;
        RECT 73.340 66.240 74.340 67.240 ;
        RECT 86.775 66.240 87.775 67.240 ;
        RECT 88.775 66.240 89.775 67.240 ;
        RECT 90.775 66.240 91.775 67.240 ;
        RECT 92.775 66.240 93.775 67.240 ;
        RECT 94.775 66.240 95.775 67.240 ;
        RECT 96.775 66.240 97.775 67.240 ;
        RECT 98.775 66.240 99.775 67.240 ;
        RECT 100.775 66.240 101.775 67.240 ;
        RECT 102.775 66.240 103.775 67.240 ;
        RECT 104.775 66.240 105.775 67.240 ;
        RECT 106.775 66.240 107.775 67.240 ;
        RECT 108.775 66.240 109.775 67.240 ;
        RECT 110.775 66.240 111.775 67.240 ;
        RECT 112.775 66.240 113.775 67.240 ;
        RECT 114.775 66.240 115.775 67.240 ;
        RECT 116.775 66.240 117.775 67.240 ;
        RECT 118.775 66.240 119.775 67.240 ;
        RECT 120.775 66.240 121.775 67.240 ;
        RECT 122.775 66.240 123.775 67.240 ;
        RECT 124.775 66.240 125.775 67.240 ;
        RECT 126.775 66.240 127.775 67.240 ;
        RECT 128.775 66.240 129.775 67.240 ;
        RECT 130.775 66.240 131.775 67.240 ;
        RECT 132.775 66.240 133.775 67.240 ;
        RECT 134.775 66.240 135.775 67.240 ;
        RECT 136.775 66.240 137.775 67.240 ;
        RECT 138.775 66.240 139.775 67.240 ;
        RECT 140.775 66.240 141.775 67.240 ;
        RECT 142.775 66.240 143.775 67.240 ;
        RECT 144.775 66.240 145.775 67.240 ;
        RECT 146.775 66.240 147.775 67.240 ;
        RECT 148.775 66.240 149.775 67.240 ;
        RECT 150.775 66.240 151.775 67.240 ;
        RECT 152.775 66.240 153.775 67.240 ;
        RECT 7.690 65.390 7.990 66.240 ;
        RECT 9.690 65.390 9.990 66.240 ;
        RECT 11.690 65.390 11.990 66.240 ;
        RECT 13.690 65.390 13.990 66.240 ;
        RECT 15.690 65.390 15.990 66.240 ;
        RECT 17.690 65.390 17.990 66.240 ;
        RECT 19.690 65.390 19.990 66.240 ;
        RECT 21.690 65.390 21.990 66.240 ;
        RECT 23.690 65.390 23.990 66.240 ;
        RECT 25.690 65.390 25.990 66.240 ;
        RECT 27.690 65.390 27.990 66.240 ;
        RECT 29.690 65.390 29.990 66.240 ;
        RECT 31.690 65.390 31.990 66.240 ;
        RECT 33.690 65.390 33.990 66.240 ;
        RECT 35.690 65.390 35.990 66.240 ;
        RECT 37.690 65.390 37.990 66.240 ;
        RECT 39.690 65.390 39.990 66.240 ;
        RECT 41.690 65.390 41.990 66.240 ;
        RECT 43.690 65.390 43.990 66.240 ;
        RECT 45.690 65.390 45.990 66.240 ;
        RECT 47.690 65.390 47.990 66.240 ;
        RECT 49.690 65.390 49.990 66.240 ;
        RECT 51.690 65.390 51.990 66.240 ;
        RECT 53.690 65.390 53.990 66.240 ;
        RECT 55.690 65.390 55.990 66.240 ;
        RECT 57.690 65.390 57.990 66.240 ;
        RECT 59.690 65.390 59.990 66.240 ;
        RECT 61.690 65.390 61.990 66.240 ;
        RECT 63.690 65.390 63.990 66.240 ;
        RECT 65.690 65.390 65.990 66.240 ;
        RECT 67.690 65.390 67.990 66.240 ;
        RECT 69.690 65.390 69.990 66.240 ;
        RECT 71.690 65.390 71.990 66.240 ;
        RECT 73.690 65.390 73.990 66.240 ;
        RECT 87.125 65.390 87.425 66.240 ;
        RECT 89.125 65.390 89.425 66.240 ;
        RECT 91.125 65.390 91.425 66.240 ;
        RECT 93.125 65.390 93.425 66.240 ;
        RECT 95.125 65.390 95.425 66.240 ;
        RECT 97.125 65.390 97.425 66.240 ;
        RECT 99.125 65.390 99.425 66.240 ;
        RECT 101.125 65.390 101.425 66.240 ;
        RECT 103.125 65.390 103.425 66.240 ;
        RECT 105.125 65.390 105.425 66.240 ;
        RECT 107.125 65.390 107.425 66.240 ;
        RECT 109.125 65.390 109.425 66.240 ;
        RECT 111.125 65.390 111.425 66.240 ;
        RECT 113.125 65.390 113.425 66.240 ;
        RECT 115.125 65.390 115.425 66.240 ;
        RECT 117.125 65.390 117.425 66.240 ;
        RECT 119.125 65.390 119.425 66.240 ;
        RECT 121.125 65.390 121.425 66.240 ;
        RECT 123.125 65.390 123.425 66.240 ;
        RECT 125.125 65.390 125.425 66.240 ;
        RECT 127.125 65.390 127.425 66.240 ;
        RECT 129.125 65.390 129.425 66.240 ;
        RECT 131.125 65.390 131.425 66.240 ;
        RECT 133.125 65.390 133.425 66.240 ;
        RECT 135.125 65.390 135.425 66.240 ;
        RECT 137.125 65.390 137.425 66.240 ;
        RECT 139.125 65.390 139.425 66.240 ;
        RECT 141.125 65.390 141.425 66.240 ;
        RECT 143.125 65.390 143.425 66.240 ;
        RECT 145.125 65.390 145.425 66.240 ;
        RECT 147.125 65.390 147.425 66.240 ;
        RECT 149.125 65.390 149.425 66.240 ;
        RECT 151.125 65.390 151.425 66.240 ;
        RECT 153.125 65.390 153.425 66.240 ;
        RECT 7.340 64.390 8.340 65.390 ;
        RECT 9.340 64.390 10.340 65.390 ;
        RECT 11.340 64.390 12.340 65.390 ;
        RECT 13.340 64.390 14.340 65.390 ;
        RECT 15.340 64.390 16.340 65.390 ;
        RECT 17.340 64.390 18.340 65.390 ;
        RECT 19.340 64.390 20.340 65.390 ;
        RECT 21.340 64.390 22.340 65.390 ;
        RECT 23.340 64.390 24.340 65.390 ;
        RECT 25.340 64.390 26.340 65.390 ;
        RECT 27.340 64.390 28.340 65.390 ;
        RECT 29.340 64.390 30.340 65.390 ;
        RECT 31.340 64.390 32.340 65.390 ;
        RECT 33.340 64.390 34.340 65.390 ;
        RECT 35.340 64.390 36.340 65.390 ;
        RECT 37.340 64.390 38.340 65.390 ;
        RECT 39.340 64.390 40.340 65.390 ;
        RECT 41.340 64.390 42.340 65.390 ;
        RECT 43.340 64.390 44.340 65.390 ;
        RECT 45.340 64.390 46.340 65.390 ;
        RECT 47.340 64.390 48.340 65.390 ;
        RECT 49.340 64.390 50.340 65.390 ;
        RECT 51.340 64.390 52.340 65.390 ;
        RECT 53.340 64.390 54.340 65.390 ;
        RECT 55.340 64.390 56.340 65.390 ;
        RECT 57.340 64.390 58.340 65.390 ;
        RECT 59.340 64.390 60.340 65.390 ;
        RECT 61.340 64.390 62.340 65.390 ;
        RECT 63.340 64.390 64.340 65.390 ;
        RECT 65.340 64.390 66.340 65.390 ;
        RECT 67.340 64.390 68.340 65.390 ;
        RECT 69.340 64.390 70.340 65.390 ;
        RECT 71.340 64.390 72.340 65.390 ;
        RECT 73.340 64.390 74.340 65.390 ;
        RECT 86.775 64.390 87.775 65.390 ;
        RECT 88.775 64.390 89.775 65.390 ;
        RECT 90.775 64.390 91.775 65.390 ;
        RECT 92.775 64.390 93.775 65.390 ;
        RECT 94.775 64.390 95.775 65.390 ;
        RECT 96.775 64.390 97.775 65.390 ;
        RECT 98.775 64.390 99.775 65.390 ;
        RECT 100.775 64.390 101.775 65.390 ;
        RECT 102.775 64.390 103.775 65.390 ;
        RECT 104.775 64.390 105.775 65.390 ;
        RECT 106.775 64.390 107.775 65.390 ;
        RECT 108.775 64.390 109.775 65.390 ;
        RECT 110.775 64.390 111.775 65.390 ;
        RECT 112.775 64.390 113.775 65.390 ;
        RECT 114.775 64.390 115.775 65.390 ;
        RECT 116.775 64.390 117.775 65.390 ;
        RECT 118.775 64.390 119.775 65.390 ;
        RECT 120.775 64.390 121.775 65.390 ;
        RECT 122.775 64.390 123.775 65.390 ;
        RECT 124.775 64.390 125.775 65.390 ;
        RECT 126.775 64.390 127.775 65.390 ;
        RECT 128.775 64.390 129.775 65.390 ;
        RECT 130.775 64.390 131.775 65.390 ;
        RECT 132.775 64.390 133.775 65.390 ;
        RECT 134.775 64.390 135.775 65.390 ;
        RECT 136.775 64.390 137.775 65.390 ;
        RECT 138.775 64.390 139.775 65.390 ;
        RECT 140.775 64.390 141.775 65.390 ;
        RECT 142.775 64.390 143.775 65.390 ;
        RECT 144.775 64.390 145.775 65.390 ;
        RECT 146.775 64.390 147.775 65.390 ;
        RECT 148.775 64.390 149.775 65.390 ;
        RECT 150.775 64.390 151.775 65.390 ;
        RECT 152.775 64.390 153.775 65.390 ;
        RECT 7.690 63.540 7.990 64.390 ;
        RECT 9.690 63.540 9.990 64.390 ;
        RECT 11.690 63.540 11.990 64.390 ;
        RECT 13.690 63.540 13.990 64.390 ;
        RECT 15.690 63.540 15.990 64.390 ;
        RECT 17.690 63.540 17.990 64.390 ;
        RECT 19.690 63.540 19.990 64.390 ;
        RECT 21.690 63.540 21.990 64.390 ;
        RECT 23.690 63.540 23.990 64.390 ;
        RECT 25.690 63.540 25.990 64.390 ;
        RECT 27.690 63.540 27.990 64.390 ;
        RECT 29.690 63.540 29.990 64.390 ;
        RECT 31.690 63.540 31.990 64.390 ;
        RECT 33.690 63.540 33.990 64.390 ;
        RECT 35.690 63.540 35.990 64.390 ;
        RECT 37.690 63.540 37.990 64.390 ;
        RECT 39.690 63.540 39.990 64.390 ;
        RECT 41.690 63.540 41.990 64.390 ;
        RECT 43.690 63.540 43.990 64.390 ;
        RECT 45.690 63.540 45.990 64.390 ;
        RECT 47.690 63.540 47.990 64.390 ;
        RECT 49.690 63.540 49.990 64.390 ;
        RECT 51.690 63.540 51.990 64.390 ;
        RECT 53.690 63.540 53.990 64.390 ;
        RECT 55.690 63.540 55.990 64.390 ;
        RECT 57.690 63.540 57.990 64.390 ;
        RECT 59.690 63.540 59.990 64.390 ;
        RECT 61.690 63.540 61.990 64.390 ;
        RECT 63.690 63.540 63.990 64.390 ;
        RECT 65.690 63.540 65.990 64.390 ;
        RECT 67.690 63.540 67.990 64.390 ;
        RECT 69.690 63.540 69.990 64.390 ;
        RECT 71.690 63.540 71.990 64.390 ;
        RECT 73.690 63.540 73.990 64.390 ;
        RECT 87.125 63.540 87.425 64.390 ;
        RECT 89.125 63.540 89.425 64.390 ;
        RECT 91.125 63.540 91.425 64.390 ;
        RECT 93.125 63.540 93.425 64.390 ;
        RECT 95.125 63.540 95.425 64.390 ;
        RECT 97.125 63.540 97.425 64.390 ;
        RECT 99.125 63.540 99.425 64.390 ;
        RECT 101.125 63.540 101.425 64.390 ;
        RECT 103.125 63.540 103.425 64.390 ;
        RECT 105.125 63.540 105.425 64.390 ;
        RECT 107.125 63.540 107.425 64.390 ;
        RECT 109.125 63.540 109.425 64.390 ;
        RECT 111.125 63.540 111.425 64.390 ;
        RECT 113.125 63.540 113.425 64.390 ;
        RECT 115.125 63.540 115.425 64.390 ;
        RECT 117.125 63.540 117.425 64.390 ;
        RECT 119.125 63.540 119.425 64.390 ;
        RECT 121.125 63.540 121.425 64.390 ;
        RECT 123.125 63.540 123.425 64.390 ;
        RECT 125.125 63.540 125.425 64.390 ;
        RECT 127.125 63.540 127.425 64.390 ;
        RECT 129.125 63.540 129.425 64.390 ;
        RECT 131.125 63.540 131.425 64.390 ;
        RECT 133.125 63.540 133.425 64.390 ;
        RECT 135.125 63.540 135.425 64.390 ;
        RECT 137.125 63.540 137.425 64.390 ;
        RECT 139.125 63.540 139.425 64.390 ;
        RECT 141.125 63.540 141.425 64.390 ;
        RECT 143.125 63.540 143.425 64.390 ;
        RECT 145.125 63.540 145.425 64.390 ;
        RECT 147.125 63.540 147.425 64.390 ;
        RECT 149.125 63.540 149.425 64.390 ;
        RECT 151.125 63.540 151.425 64.390 ;
        RECT 153.125 63.540 153.425 64.390 ;
        RECT 7.340 62.540 8.340 63.540 ;
        RECT 9.340 62.540 10.340 63.540 ;
        RECT 11.340 62.540 12.340 63.540 ;
        RECT 13.340 62.540 14.340 63.540 ;
        RECT 15.340 62.540 16.340 63.540 ;
        RECT 17.340 62.540 18.340 63.540 ;
        RECT 19.340 62.540 20.340 63.540 ;
        RECT 21.340 62.540 22.340 63.540 ;
        RECT 23.340 62.540 24.340 63.540 ;
        RECT 25.340 62.540 26.340 63.540 ;
        RECT 27.340 62.540 28.340 63.540 ;
        RECT 29.340 62.540 30.340 63.540 ;
        RECT 31.340 62.540 32.340 63.540 ;
        RECT 33.340 62.540 34.340 63.540 ;
        RECT 35.340 62.540 36.340 63.540 ;
        RECT 37.340 62.540 38.340 63.540 ;
        RECT 39.340 62.540 40.340 63.540 ;
        RECT 41.340 62.540 42.340 63.540 ;
        RECT 43.340 62.540 44.340 63.540 ;
        RECT 45.340 62.540 46.340 63.540 ;
        RECT 47.340 62.540 48.340 63.540 ;
        RECT 49.340 62.540 50.340 63.540 ;
        RECT 51.340 62.540 52.340 63.540 ;
        RECT 53.340 62.540 54.340 63.540 ;
        RECT 55.340 62.540 56.340 63.540 ;
        RECT 57.340 62.540 58.340 63.540 ;
        RECT 59.340 62.540 60.340 63.540 ;
        RECT 61.340 62.540 62.340 63.540 ;
        RECT 63.340 62.540 64.340 63.540 ;
        RECT 65.340 62.540 66.340 63.540 ;
        RECT 67.340 62.540 68.340 63.540 ;
        RECT 69.340 62.540 70.340 63.540 ;
        RECT 71.340 62.540 72.340 63.540 ;
        RECT 73.340 62.540 74.340 63.540 ;
        RECT 86.775 62.540 87.775 63.540 ;
        RECT 88.775 62.540 89.775 63.540 ;
        RECT 90.775 62.540 91.775 63.540 ;
        RECT 92.775 62.540 93.775 63.540 ;
        RECT 94.775 62.540 95.775 63.540 ;
        RECT 96.775 62.540 97.775 63.540 ;
        RECT 98.775 62.540 99.775 63.540 ;
        RECT 100.775 62.540 101.775 63.540 ;
        RECT 102.775 62.540 103.775 63.540 ;
        RECT 104.775 62.540 105.775 63.540 ;
        RECT 106.775 62.540 107.775 63.540 ;
        RECT 108.775 62.540 109.775 63.540 ;
        RECT 110.775 62.540 111.775 63.540 ;
        RECT 112.775 62.540 113.775 63.540 ;
        RECT 114.775 62.540 115.775 63.540 ;
        RECT 116.775 62.540 117.775 63.540 ;
        RECT 118.775 62.540 119.775 63.540 ;
        RECT 120.775 62.540 121.775 63.540 ;
        RECT 122.775 62.540 123.775 63.540 ;
        RECT 124.775 62.540 125.775 63.540 ;
        RECT 126.775 62.540 127.775 63.540 ;
        RECT 128.775 62.540 129.775 63.540 ;
        RECT 130.775 62.540 131.775 63.540 ;
        RECT 132.775 62.540 133.775 63.540 ;
        RECT 134.775 62.540 135.775 63.540 ;
        RECT 136.775 62.540 137.775 63.540 ;
        RECT 138.775 62.540 139.775 63.540 ;
        RECT 140.775 62.540 141.775 63.540 ;
        RECT 142.775 62.540 143.775 63.540 ;
        RECT 144.775 62.540 145.775 63.540 ;
        RECT 146.775 62.540 147.775 63.540 ;
        RECT 148.775 62.540 149.775 63.540 ;
        RECT 150.775 62.540 151.775 63.540 ;
        RECT 152.775 62.540 153.775 63.540 ;
        RECT 7.690 61.690 7.990 62.540 ;
        RECT 9.690 61.690 9.990 62.540 ;
        RECT 11.690 61.690 11.990 62.540 ;
        RECT 13.690 61.690 13.990 62.540 ;
        RECT 15.690 61.690 15.990 62.540 ;
        RECT 17.690 61.690 17.990 62.540 ;
        RECT 19.690 61.690 19.990 62.540 ;
        RECT 21.690 61.690 21.990 62.540 ;
        RECT 23.690 61.690 23.990 62.540 ;
        RECT 25.690 61.690 25.990 62.540 ;
        RECT 27.690 61.690 27.990 62.540 ;
        RECT 29.690 61.690 29.990 62.540 ;
        RECT 31.690 61.690 31.990 62.540 ;
        RECT 33.690 61.690 33.990 62.540 ;
        RECT 35.690 61.690 35.990 62.540 ;
        RECT 37.690 61.690 37.990 62.540 ;
        RECT 39.690 61.690 39.990 62.540 ;
        RECT 41.690 61.690 41.990 62.540 ;
        RECT 43.690 61.690 43.990 62.540 ;
        RECT 45.690 61.690 45.990 62.540 ;
        RECT 47.690 61.690 47.990 62.540 ;
        RECT 49.690 61.690 49.990 62.540 ;
        RECT 51.690 61.690 51.990 62.540 ;
        RECT 53.690 61.690 53.990 62.540 ;
        RECT 55.690 61.690 55.990 62.540 ;
        RECT 57.690 61.690 57.990 62.540 ;
        RECT 59.690 61.690 59.990 62.540 ;
        RECT 61.690 61.690 61.990 62.540 ;
        RECT 63.690 61.690 63.990 62.540 ;
        RECT 65.690 61.690 65.990 62.540 ;
        RECT 67.690 61.690 67.990 62.540 ;
        RECT 69.690 61.690 69.990 62.540 ;
        RECT 71.690 61.690 71.990 62.540 ;
        RECT 73.690 61.690 73.990 62.540 ;
        RECT 87.125 61.690 87.425 62.540 ;
        RECT 89.125 61.690 89.425 62.540 ;
        RECT 91.125 61.690 91.425 62.540 ;
        RECT 93.125 61.690 93.425 62.540 ;
        RECT 95.125 61.690 95.425 62.540 ;
        RECT 97.125 61.690 97.425 62.540 ;
        RECT 99.125 61.690 99.425 62.540 ;
        RECT 101.125 61.690 101.425 62.540 ;
        RECT 103.125 61.690 103.425 62.540 ;
        RECT 105.125 61.690 105.425 62.540 ;
        RECT 107.125 61.690 107.425 62.540 ;
        RECT 109.125 61.690 109.425 62.540 ;
        RECT 111.125 61.690 111.425 62.540 ;
        RECT 113.125 61.690 113.425 62.540 ;
        RECT 115.125 61.690 115.425 62.540 ;
        RECT 117.125 61.690 117.425 62.540 ;
        RECT 119.125 61.690 119.425 62.540 ;
        RECT 121.125 61.690 121.425 62.540 ;
        RECT 123.125 61.690 123.425 62.540 ;
        RECT 125.125 61.690 125.425 62.540 ;
        RECT 127.125 61.690 127.425 62.540 ;
        RECT 129.125 61.690 129.425 62.540 ;
        RECT 131.125 61.690 131.425 62.540 ;
        RECT 133.125 61.690 133.425 62.540 ;
        RECT 135.125 61.690 135.425 62.540 ;
        RECT 137.125 61.690 137.425 62.540 ;
        RECT 139.125 61.690 139.425 62.540 ;
        RECT 141.125 61.690 141.425 62.540 ;
        RECT 143.125 61.690 143.425 62.540 ;
        RECT 145.125 61.690 145.425 62.540 ;
        RECT 147.125 61.690 147.425 62.540 ;
        RECT 149.125 61.690 149.425 62.540 ;
        RECT 151.125 61.690 151.425 62.540 ;
        RECT 153.125 61.690 153.425 62.540 ;
        RECT 7.340 60.690 8.340 61.690 ;
        RECT 9.340 60.690 10.340 61.690 ;
        RECT 11.340 60.690 12.340 61.690 ;
        RECT 13.340 60.690 14.340 61.690 ;
        RECT 15.340 60.690 16.340 61.690 ;
        RECT 17.340 60.690 18.340 61.690 ;
        RECT 19.340 60.690 20.340 61.690 ;
        RECT 21.340 60.690 22.340 61.690 ;
        RECT 23.340 60.690 24.340 61.690 ;
        RECT 25.340 60.690 26.340 61.690 ;
        RECT 27.340 60.690 28.340 61.690 ;
        RECT 29.340 60.690 30.340 61.690 ;
        RECT 31.340 60.690 32.340 61.690 ;
        RECT 33.340 60.690 34.340 61.690 ;
        RECT 35.340 60.690 36.340 61.690 ;
        RECT 37.340 60.690 38.340 61.690 ;
        RECT 39.340 60.690 40.340 61.690 ;
        RECT 41.340 60.690 42.340 61.690 ;
        RECT 43.340 60.690 44.340 61.690 ;
        RECT 45.340 60.690 46.340 61.690 ;
        RECT 47.340 60.690 48.340 61.690 ;
        RECT 49.340 60.690 50.340 61.690 ;
        RECT 51.340 60.690 52.340 61.690 ;
        RECT 53.340 60.690 54.340 61.690 ;
        RECT 55.340 60.690 56.340 61.690 ;
        RECT 57.340 60.690 58.340 61.690 ;
        RECT 59.340 60.690 60.340 61.690 ;
        RECT 61.340 60.690 62.340 61.690 ;
        RECT 63.340 60.690 64.340 61.690 ;
        RECT 65.340 60.690 66.340 61.690 ;
        RECT 67.340 60.690 68.340 61.690 ;
        RECT 69.340 60.690 70.340 61.690 ;
        RECT 71.340 60.690 72.340 61.690 ;
        RECT 73.340 60.690 74.340 61.690 ;
        RECT 86.775 60.690 87.775 61.690 ;
        RECT 88.775 60.690 89.775 61.690 ;
        RECT 90.775 60.690 91.775 61.690 ;
        RECT 92.775 60.690 93.775 61.690 ;
        RECT 94.775 60.690 95.775 61.690 ;
        RECT 96.775 60.690 97.775 61.690 ;
        RECT 98.775 60.690 99.775 61.690 ;
        RECT 100.775 60.690 101.775 61.690 ;
        RECT 102.775 60.690 103.775 61.690 ;
        RECT 104.775 60.690 105.775 61.690 ;
        RECT 106.775 60.690 107.775 61.690 ;
        RECT 108.775 60.690 109.775 61.690 ;
        RECT 110.775 60.690 111.775 61.690 ;
        RECT 112.775 60.690 113.775 61.690 ;
        RECT 114.775 60.690 115.775 61.690 ;
        RECT 116.775 60.690 117.775 61.690 ;
        RECT 118.775 60.690 119.775 61.690 ;
        RECT 120.775 60.690 121.775 61.690 ;
        RECT 122.775 60.690 123.775 61.690 ;
        RECT 124.775 60.690 125.775 61.690 ;
        RECT 126.775 60.690 127.775 61.690 ;
        RECT 128.775 60.690 129.775 61.690 ;
        RECT 130.775 60.690 131.775 61.690 ;
        RECT 132.775 60.690 133.775 61.690 ;
        RECT 134.775 60.690 135.775 61.690 ;
        RECT 136.775 60.690 137.775 61.690 ;
        RECT 138.775 60.690 139.775 61.690 ;
        RECT 140.775 60.690 141.775 61.690 ;
        RECT 142.775 60.690 143.775 61.690 ;
        RECT 144.775 60.690 145.775 61.690 ;
        RECT 146.775 60.690 147.775 61.690 ;
        RECT 148.775 60.690 149.775 61.690 ;
        RECT 150.775 60.690 151.775 61.690 ;
        RECT 152.775 60.690 153.775 61.690 ;
        RECT 7.690 59.840 7.990 60.690 ;
        RECT 9.690 59.840 9.990 60.690 ;
        RECT 11.690 59.840 11.990 60.690 ;
        RECT 13.690 59.840 13.990 60.690 ;
        RECT 15.690 59.840 15.990 60.690 ;
        RECT 17.690 59.840 17.990 60.690 ;
        RECT 19.690 59.840 19.990 60.690 ;
        RECT 21.690 59.840 21.990 60.690 ;
        RECT 23.690 59.840 23.990 60.690 ;
        RECT 25.690 59.840 25.990 60.690 ;
        RECT 27.690 59.840 27.990 60.690 ;
        RECT 29.690 59.840 29.990 60.690 ;
        RECT 31.690 59.840 31.990 60.690 ;
        RECT 33.690 59.840 33.990 60.690 ;
        RECT 35.690 59.840 35.990 60.690 ;
        RECT 37.690 59.840 37.990 60.690 ;
        RECT 39.690 59.840 39.990 60.690 ;
        RECT 41.690 59.840 41.990 60.690 ;
        RECT 43.690 59.840 43.990 60.690 ;
        RECT 45.690 59.840 45.990 60.690 ;
        RECT 47.690 59.840 47.990 60.690 ;
        RECT 49.690 59.840 49.990 60.690 ;
        RECT 51.690 59.840 51.990 60.690 ;
        RECT 53.690 59.840 53.990 60.690 ;
        RECT 55.690 59.840 55.990 60.690 ;
        RECT 57.690 59.840 57.990 60.690 ;
        RECT 59.690 59.840 59.990 60.690 ;
        RECT 61.690 59.840 61.990 60.690 ;
        RECT 63.690 59.840 63.990 60.690 ;
        RECT 65.690 59.840 65.990 60.690 ;
        RECT 67.690 59.840 67.990 60.690 ;
        RECT 69.690 59.840 69.990 60.690 ;
        RECT 71.690 59.840 71.990 60.690 ;
        RECT 73.690 59.840 73.990 60.690 ;
        RECT 87.125 59.840 87.425 60.690 ;
        RECT 89.125 59.840 89.425 60.690 ;
        RECT 91.125 59.840 91.425 60.690 ;
        RECT 93.125 59.840 93.425 60.690 ;
        RECT 95.125 59.840 95.425 60.690 ;
        RECT 97.125 59.840 97.425 60.690 ;
        RECT 99.125 59.840 99.425 60.690 ;
        RECT 101.125 59.840 101.425 60.690 ;
        RECT 103.125 59.840 103.425 60.690 ;
        RECT 105.125 59.840 105.425 60.690 ;
        RECT 107.125 59.840 107.425 60.690 ;
        RECT 109.125 59.840 109.425 60.690 ;
        RECT 111.125 59.840 111.425 60.690 ;
        RECT 113.125 59.840 113.425 60.690 ;
        RECT 115.125 59.840 115.425 60.690 ;
        RECT 117.125 59.840 117.425 60.690 ;
        RECT 119.125 59.840 119.425 60.690 ;
        RECT 121.125 59.840 121.425 60.690 ;
        RECT 123.125 59.840 123.425 60.690 ;
        RECT 125.125 59.840 125.425 60.690 ;
        RECT 127.125 59.840 127.425 60.690 ;
        RECT 129.125 59.840 129.425 60.690 ;
        RECT 131.125 59.840 131.425 60.690 ;
        RECT 133.125 59.840 133.425 60.690 ;
        RECT 135.125 59.840 135.425 60.690 ;
        RECT 137.125 59.840 137.425 60.690 ;
        RECT 139.125 59.840 139.425 60.690 ;
        RECT 141.125 59.840 141.425 60.690 ;
        RECT 143.125 59.840 143.425 60.690 ;
        RECT 145.125 59.840 145.425 60.690 ;
        RECT 147.125 59.840 147.425 60.690 ;
        RECT 149.125 59.840 149.425 60.690 ;
        RECT 151.125 59.840 151.425 60.690 ;
        RECT 153.125 59.840 153.425 60.690 ;
        RECT 7.340 58.840 8.340 59.840 ;
        RECT 9.340 58.840 10.340 59.840 ;
        RECT 11.340 58.840 12.340 59.840 ;
        RECT 13.340 58.840 14.340 59.840 ;
        RECT 15.340 58.840 16.340 59.840 ;
        RECT 17.340 58.840 18.340 59.840 ;
        RECT 19.340 58.840 20.340 59.840 ;
        RECT 21.340 58.840 22.340 59.840 ;
        RECT 23.340 58.840 24.340 59.840 ;
        RECT 25.340 58.840 26.340 59.840 ;
        RECT 27.340 58.840 28.340 59.840 ;
        RECT 29.340 58.840 30.340 59.840 ;
        RECT 31.340 58.840 32.340 59.840 ;
        RECT 33.340 58.840 34.340 59.840 ;
        RECT 35.340 58.840 36.340 59.840 ;
        RECT 37.340 58.840 38.340 59.840 ;
        RECT 39.340 58.840 40.340 59.840 ;
        RECT 41.340 58.840 42.340 59.840 ;
        RECT 43.340 58.840 44.340 59.840 ;
        RECT 45.340 58.840 46.340 59.840 ;
        RECT 47.340 58.840 48.340 59.840 ;
        RECT 49.340 58.840 50.340 59.840 ;
        RECT 51.340 58.840 52.340 59.840 ;
        RECT 53.340 58.840 54.340 59.840 ;
        RECT 55.340 58.840 56.340 59.840 ;
        RECT 57.340 58.840 58.340 59.840 ;
        RECT 59.340 58.840 60.340 59.840 ;
        RECT 61.340 58.840 62.340 59.840 ;
        RECT 63.340 58.840 64.340 59.840 ;
        RECT 65.340 58.840 66.340 59.840 ;
        RECT 67.340 58.840 68.340 59.840 ;
        RECT 69.340 58.840 70.340 59.840 ;
        RECT 71.340 58.840 72.340 59.840 ;
        RECT 73.340 58.840 74.340 59.840 ;
        RECT 86.775 58.840 87.775 59.840 ;
        RECT 88.775 58.840 89.775 59.840 ;
        RECT 90.775 58.840 91.775 59.840 ;
        RECT 92.775 58.840 93.775 59.840 ;
        RECT 94.775 58.840 95.775 59.840 ;
        RECT 96.775 58.840 97.775 59.840 ;
        RECT 98.775 58.840 99.775 59.840 ;
        RECT 100.775 58.840 101.775 59.840 ;
        RECT 102.775 58.840 103.775 59.840 ;
        RECT 104.775 58.840 105.775 59.840 ;
        RECT 106.775 58.840 107.775 59.840 ;
        RECT 108.775 58.840 109.775 59.840 ;
        RECT 110.775 58.840 111.775 59.840 ;
        RECT 112.775 58.840 113.775 59.840 ;
        RECT 114.775 58.840 115.775 59.840 ;
        RECT 116.775 58.840 117.775 59.840 ;
        RECT 118.775 58.840 119.775 59.840 ;
        RECT 120.775 58.840 121.775 59.840 ;
        RECT 122.775 58.840 123.775 59.840 ;
        RECT 124.775 58.840 125.775 59.840 ;
        RECT 126.775 58.840 127.775 59.840 ;
        RECT 128.775 58.840 129.775 59.840 ;
        RECT 130.775 58.840 131.775 59.840 ;
        RECT 132.775 58.840 133.775 59.840 ;
        RECT 134.775 58.840 135.775 59.840 ;
        RECT 136.775 58.840 137.775 59.840 ;
        RECT 138.775 58.840 139.775 59.840 ;
        RECT 140.775 58.840 141.775 59.840 ;
        RECT 142.775 58.840 143.775 59.840 ;
        RECT 144.775 58.840 145.775 59.840 ;
        RECT 146.775 58.840 147.775 59.840 ;
        RECT 148.775 58.840 149.775 59.840 ;
        RECT 150.775 58.840 151.775 59.840 ;
        RECT 152.775 58.840 153.775 59.840 ;
        RECT 7.690 57.990 7.990 58.840 ;
        RECT 9.690 57.990 9.990 58.840 ;
        RECT 11.690 57.990 11.990 58.840 ;
        RECT 13.690 57.990 13.990 58.840 ;
        RECT 15.690 57.990 15.990 58.840 ;
        RECT 17.690 57.990 17.990 58.840 ;
        RECT 19.690 57.990 19.990 58.840 ;
        RECT 21.690 57.990 21.990 58.840 ;
        RECT 23.690 57.990 23.990 58.840 ;
        RECT 25.690 57.990 25.990 58.840 ;
        RECT 27.690 57.990 27.990 58.840 ;
        RECT 29.690 57.990 29.990 58.840 ;
        RECT 31.690 57.990 31.990 58.840 ;
        RECT 33.690 57.990 33.990 58.840 ;
        RECT 35.690 57.990 35.990 58.840 ;
        RECT 37.690 57.990 37.990 58.840 ;
        RECT 39.690 57.990 39.990 58.840 ;
        RECT 41.690 57.990 41.990 58.840 ;
        RECT 43.690 57.990 43.990 58.840 ;
        RECT 45.690 57.990 45.990 58.840 ;
        RECT 47.690 57.990 47.990 58.840 ;
        RECT 49.690 57.990 49.990 58.840 ;
        RECT 51.690 57.990 51.990 58.840 ;
        RECT 53.690 57.990 53.990 58.840 ;
        RECT 55.690 57.990 55.990 58.840 ;
        RECT 57.690 57.990 57.990 58.840 ;
        RECT 59.690 57.990 59.990 58.840 ;
        RECT 61.690 57.990 61.990 58.840 ;
        RECT 63.690 57.990 63.990 58.840 ;
        RECT 65.690 57.990 65.990 58.840 ;
        RECT 67.690 57.990 67.990 58.840 ;
        RECT 69.690 57.990 69.990 58.840 ;
        RECT 71.690 57.990 71.990 58.840 ;
        RECT 73.690 57.990 73.990 58.840 ;
        RECT 87.125 57.990 87.425 58.840 ;
        RECT 89.125 57.990 89.425 58.840 ;
        RECT 91.125 57.990 91.425 58.840 ;
        RECT 93.125 57.990 93.425 58.840 ;
        RECT 95.125 57.990 95.425 58.840 ;
        RECT 97.125 57.990 97.425 58.840 ;
        RECT 99.125 57.990 99.425 58.840 ;
        RECT 101.125 57.990 101.425 58.840 ;
        RECT 103.125 57.990 103.425 58.840 ;
        RECT 105.125 57.990 105.425 58.840 ;
        RECT 107.125 57.990 107.425 58.840 ;
        RECT 109.125 57.990 109.425 58.840 ;
        RECT 111.125 57.990 111.425 58.840 ;
        RECT 113.125 57.990 113.425 58.840 ;
        RECT 115.125 57.990 115.425 58.840 ;
        RECT 117.125 57.990 117.425 58.840 ;
        RECT 119.125 57.990 119.425 58.840 ;
        RECT 121.125 57.990 121.425 58.840 ;
        RECT 123.125 57.990 123.425 58.840 ;
        RECT 125.125 57.990 125.425 58.840 ;
        RECT 127.125 57.990 127.425 58.840 ;
        RECT 129.125 57.990 129.425 58.840 ;
        RECT 131.125 57.990 131.425 58.840 ;
        RECT 133.125 57.990 133.425 58.840 ;
        RECT 135.125 57.990 135.425 58.840 ;
        RECT 137.125 57.990 137.425 58.840 ;
        RECT 139.125 57.990 139.425 58.840 ;
        RECT 141.125 57.990 141.425 58.840 ;
        RECT 143.125 57.990 143.425 58.840 ;
        RECT 145.125 57.990 145.425 58.840 ;
        RECT 147.125 57.990 147.425 58.840 ;
        RECT 149.125 57.990 149.425 58.840 ;
        RECT 151.125 57.990 151.425 58.840 ;
        RECT 153.125 57.990 153.425 58.840 ;
        RECT 7.340 56.990 8.340 57.990 ;
        RECT 9.340 56.990 10.340 57.990 ;
        RECT 11.340 56.990 12.340 57.990 ;
        RECT 13.340 56.990 14.340 57.990 ;
        RECT 15.340 56.990 16.340 57.990 ;
        RECT 17.340 56.990 18.340 57.990 ;
        RECT 19.340 56.990 20.340 57.990 ;
        RECT 21.340 56.990 22.340 57.990 ;
        RECT 23.340 56.990 24.340 57.990 ;
        RECT 25.340 56.990 26.340 57.990 ;
        RECT 27.340 56.990 28.340 57.990 ;
        RECT 29.340 56.990 30.340 57.990 ;
        RECT 31.340 56.990 32.340 57.990 ;
        RECT 33.340 56.990 34.340 57.990 ;
        RECT 35.340 56.990 36.340 57.990 ;
        RECT 37.340 56.990 38.340 57.990 ;
        RECT 39.340 56.990 40.340 57.990 ;
        RECT 41.340 56.990 42.340 57.990 ;
        RECT 43.340 56.990 44.340 57.990 ;
        RECT 45.340 56.990 46.340 57.990 ;
        RECT 47.340 56.990 48.340 57.990 ;
        RECT 49.340 56.990 50.340 57.990 ;
        RECT 51.340 56.990 52.340 57.990 ;
        RECT 53.340 56.990 54.340 57.990 ;
        RECT 55.340 56.990 56.340 57.990 ;
        RECT 57.340 56.990 58.340 57.990 ;
        RECT 59.340 56.990 60.340 57.990 ;
        RECT 61.340 56.990 62.340 57.990 ;
        RECT 63.340 56.990 64.340 57.990 ;
        RECT 65.340 56.990 66.340 57.990 ;
        RECT 67.340 56.990 68.340 57.990 ;
        RECT 69.340 56.990 70.340 57.990 ;
        RECT 71.340 56.990 72.340 57.990 ;
        RECT 73.340 56.990 74.340 57.990 ;
        RECT 86.775 56.990 87.775 57.990 ;
        RECT 88.775 56.990 89.775 57.990 ;
        RECT 90.775 56.990 91.775 57.990 ;
        RECT 92.775 56.990 93.775 57.990 ;
        RECT 94.775 56.990 95.775 57.990 ;
        RECT 96.775 56.990 97.775 57.990 ;
        RECT 98.775 56.990 99.775 57.990 ;
        RECT 100.775 56.990 101.775 57.990 ;
        RECT 102.775 56.990 103.775 57.990 ;
        RECT 104.775 56.990 105.775 57.990 ;
        RECT 106.775 56.990 107.775 57.990 ;
        RECT 108.775 56.990 109.775 57.990 ;
        RECT 110.775 56.990 111.775 57.990 ;
        RECT 112.775 56.990 113.775 57.990 ;
        RECT 114.775 56.990 115.775 57.990 ;
        RECT 116.775 56.990 117.775 57.990 ;
        RECT 118.775 56.990 119.775 57.990 ;
        RECT 120.775 56.990 121.775 57.990 ;
        RECT 122.775 56.990 123.775 57.990 ;
        RECT 124.775 56.990 125.775 57.990 ;
        RECT 126.775 56.990 127.775 57.990 ;
        RECT 128.775 56.990 129.775 57.990 ;
        RECT 130.775 56.990 131.775 57.990 ;
        RECT 132.775 56.990 133.775 57.990 ;
        RECT 134.775 56.990 135.775 57.990 ;
        RECT 136.775 56.990 137.775 57.990 ;
        RECT 138.775 56.990 139.775 57.990 ;
        RECT 140.775 56.990 141.775 57.990 ;
        RECT 142.775 56.990 143.775 57.990 ;
        RECT 144.775 56.990 145.775 57.990 ;
        RECT 146.775 56.990 147.775 57.990 ;
        RECT 148.775 56.990 149.775 57.990 ;
        RECT 150.775 56.990 151.775 57.990 ;
        RECT 152.775 56.990 153.775 57.990 ;
        RECT 7.690 56.140 7.990 56.990 ;
        RECT 9.690 56.140 9.990 56.990 ;
        RECT 11.690 56.140 11.990 56.990 ;
        RECT 13.690 56.140 13.990 56.990 ;
        RECT 15.690 56.140 15.990 56.990 ;
        RECT 17.690 56.140 17.990 56.990 ;
        RECT 19.690 56.140 19.990 56.990 ;
        RECT 21.690 56.140 21.990 56.990 ;
        RECT 23.690 56.140 23.990 56.990 ;
        RECT 25.690 56.140 25.990 56.990 ;
        RECT 27.690 56.140 27.990 56.990 ;
        RECT 29.690 56.140 29.990 56.990 ;
        RECT 31.690 56.140 31.990 56.990 ;
        RECT 33.690 56.140 33.990 56.990 ;
        RECT 35.690 56.140 35.990 56.990 ;
        RECT 37.690 56.140 37.990 56.990 ;
        RECT 39.690 56.140 39.990 56.990 ;
        RECT 41.690 56.140 41.990 56.990 ;
        RECT 43.690 56.140 43.990 56.990 ;
        RECT 45.690 56.140 45.990 56.990 ;
        RECT 47.690 56.140 47.990 56.990 ;
        RECT 49.690 56.140 49.990 56.990 ;
        RECT 51.690 56.140 51.990 56.990 ;
        RECT 53.690 56.140 53.990 56.990 ;
        RECT 55.690 56.140 55.990 56.990 ;
        RECT 57.690 56.140 57.990 56.990 ;
        RECT 59.690 56.140 59.990 56.990 ;
        RECT 61.690 56.140 61.990 56.990 ;
        RECT 63.690 56.140 63.990 56.990 ;
        RECT 65.690 56.140 65.990 56.990 ;
        RECT 67.690 56.140 67.990 56.990 ;
        RECT 69.690 56.140 69.990 56.990 ;
        RECT 71.690 56.140 71.990 56.990 ;
        RECT 73.690 56.140 73.990 56.990 ;
        RECT 87.125 56.140 87.425 56.990 ;
        RECT 89.125 56.140 89.425 56.990 ;
        RECT 91.125 56.140 91.425 56.990 ;
        RECT 93.125 56.140 93.425 56.990 ;
        RECT 95.125 56.140 95.425 56.990 ;
        RECT 97.125 56.140 97.425 56.990 ;
        RECT 99.125 56.140 99.425 56.990 ;
        RECT 101.125 56.140 101.425 56.990 ;
        RECT 103.125 56.140 103.425 56.990 ;
        RECT 105.125 56.140 105.425 56.990 ;
        RECT 107.125 56.140 107.425 56.990 ;
        RECT 109.125 56.140 109.425 56.990 ;
        RECT 111.125 56.140 111.425 56.990 ;
        RECT 113.125 56.140 113.425 56.990 ;
        RECT 115.125 56.140 115.425 56.990 ;
        RECT 117.125 56.140 117.425 56.990 ;
        RECT 119.125 56.140 119.425 56.990 ;
        RECT 121.125 56.140 121.425 56.990 ;
        RECT 123.125 56.140 123.425 56.990 ;
        RECT 125.125 56.140 125.425 56.990 ;
        RECT 127.125 56.140 127.425 56.990 ;
        RECT 129.125 56.140 129.425 56.990 ;
        RECT 131.125 56.140 131.425 56.990 ;
        RECT 133.125 56.140 133.425 56.990 ;
        RECT 135.125 56.140 135.425 56.990 ;
        RECT 137.125 56.140 137.425 56.990 ;
        RECT 139.125 56.140 139.425 56.990 ;
        RECT 141.125 56.140 141.425 56.990 ;
        RECT 143.125 56.140 143.425 56.990 ;
        RECT 145.125 56.140 145.425 56.990 ;
        RECT 147.125 56.140 147.425 56.990 ;
        RECT 149.125 56.140 149.425 56.990 ;
        RECT 151.125 56.140 151.425 56.990 ;
        RECT 153.125 56.140 153.425 56.990 ;
        RECT 7.340 55.140 8.340 56.140 ;
        RECT 9.340 55.140 10.340 56.140 ;
        RECT 11.340 55.140 12.340 56.140 ;
        RECT 13.340 55.140 14.340 56.140 ;
        RECT 15.340 55.140 16.340 56.140 ;
        RECT 17.340 55.140 18.340 56.140 ;
        RECT 19.340 55.140 20.340 56.140 ;
        RECT 21.340 55.140 22.340 56.140 ;
        RECT 23.340 55.140 24.340 56.140 ;
        RECT 25.340 55.140 26.340 56.140 ;
        RECT 27.340 55.140 28.340 56.140 ;
        RECT 29.340 55.140 30.340 56.140 ;
        RECT 31.340 55.140 32.340 56.140 ;
        RECT 33.340 55.140 34.340 56.140 ;
        RECT 35.340 55.140 36.340 56.140 ;
        RECT 37.340 55.140 38.340 56.140 ;
        RECT 39.340 55.140 40.340 56.140 ;
        RECT 41.340 55.140 42.340 56.140 ;
        RECT 43.340 55.140 44.340 56.140 ;
        RECT 45.340 55.140 46.340 56.140 ;
        RECT 47.340 55.140 48.340 56.140 ;
        RECT 49.340 55.140 50.340 56.140 ;
        RECT 51.340 55.140 52.340 56.140 ;
        RECT 53.340 55.140 54.340 56.140 ;
        RECT 55.340 55.140 56.340 56.140 ;
        RECT 57.340 55.140 58.340 56.140 ;
        RECT 59.340 55.140 60.340 56.140 ;
        RECT 61.340 55.140 62.340 56.140 ;
        RECT 63.340 55.140 64.340 56.140 ;
        RECT 65.340 55.140 66.340 56.140 ;
        RECT 67.340 55.140 68.340 56.140 ;
        RECT 69.340 55.140 70.340 56.140 ;
        RECT 71.340 55.140 72.340 56.140 ;
        RECT 73.340 55.140 74.340 56.140 ;
        RECT 86.775 55.140 87.775 56.140 ;
        RECT 88.775 55.140 89.775 56.140 ;
        RECT 90.775 55.140 91.775 56.140 ;
        RECT 92.775 55.140 93.775 56.140 ;
        RECT 94.775 55.140 95.775 56.140 ;
        RECT 96.775 55.140 97.775 56.140 ;
        RECT 98.775 55.140 99.775 56.140 ;
        RECT 100.775 55.140 101.775 56.140 ;
        RECT 102.775 55.140 103.775 56.140 ;
        RECT 104.775 55.140 105.775 56.140 ;
        RECT 106.775 55.140 107.775 56.140 ;
        RECT 108.775 55.140 109.775 56.140 ;
        RECT 110.775 55.140 111.775 56.140 ;
        RECT 112.775 55.140 113.775 56.140 ;
        RECT 114.775 55.140 115.775 56.140 ;
        RECT 116.775 55.140 117.775 56.140 ;
        RECT 118.775 55.140 119.775 56.140 ;
        RECT 120.775 55.140 121.775 56.140 ;
        RECT 122.775 55.140 123.775 56.140 ;
        RECT 124.775 55.140 125.775 56.140 ;
        RECT 126.775 55.140 127.775 56.140 ;
        RECT 128.775 55.140 129.775 56.140 ;
        RECT 130.775 55.140 131.775 56.140 ;
        RECT 132.775 55.140 133.775 56.140 ;
        RECT 134.775 55.140 135.775 56.140 ;
        RECT 136.775 55.140 137.775 56.140 ;
        RECT 138.775 55.140 139.775 56.140 ;
        RECT 140.775 55.140 141.775 56.140 ;
        RECT 142.775 55.140 143.775 56.140 ;
        RECT 144.775 55.140 145.775 56.140 ;
        RECT 146.775 55.140 147.775 56.140 ;
        RECT 148.775 55.140 149.775 56.140 ;
        RECT 150.775 55.140 151.775 56.140 ;
        RECT 152.775 55.140 153.775 56.140 ;
        RECT 7.690 54.290 7.990 55.140 ;
        RECT 9.690 54.290 9.990 55.140 ;
        RECT 11.690 54.290 11.990 55.140 ;
        RECT 13.690 54.290 13.990 55.140 ;
        RECT 15.690 54.290 15.990 55.140 ;
        RECT 17.690 54.290 17.990 55.140 ;
        RECT 19.690 54.290 19.990 55.140 ;
        RECT 21.690 54.290 21.990 55.140 ;
        RECT 23.690 54.290 23.990 55.140 ;
        RECT 25.690 54.290 25.990 55.140 ;
        RECT 27.690 54.290 27.990 55.140 ;
        RECT 29.690 54.290 29.990 55.140 ;
        RECT 31.690 54.290 31.990 55.140 ;
        RECT 33.690 54.290 33.990 55.140 ;
        RECT 35.690 54.290 35.990 55.140 ;
        RECT 37.690 54.290 37.990 55.140 ;
        RECT 39.690 54.290 39.990 55.140 ;
        RECT 41.690 54.290 41.990 55.140 ;
        RECT 43.690 54.290 43.990 55.140 ;
        RECT 45.690 54.290 45.990 55.140 ;
        RECT 47.690 54.290 47.990 55.140 ;
        RECT 49.690 54.290 49.990 55.140 ;
        RECT 51.690 54.290 51.990 55.140 ;
        RECT 53.690 54.290 53.990 55.140 ;
        RECT 55.690 54.290 55.990 55.140 ;
        RECT 57.690 54.290 57.990 55.140 ;
        RECT 59.690 54.290 59.990 55.140 ;
        RECT 61.690 54.290 61.990 55.140 ;
        RECT 63.690 54.290 63.990 55.140 ;
        RECT 65.690 54.290 65.990 55.140 ;
        RECT 67.690 54.290 67.990 55.140 ;
        RECT 69.690 54.290 69.990 55.140 ;
        RECT 71.690 54.290 71.990 55.140 ;
        RECT 73.690 54.290 73.990 55.140 ;
        RECT 87.125 54.290 87.425 55.140 ;
        RECT 89.125 54.290 89.425 55.140 ;
        RECT 91.125 54.290 91.425 55.140 ;
        RECT 93.125 54.290 93.425 55.140 ;
        RECT 95.125 54.290 95.425 55.140 ;
        RECT 97.125 54.290 97.425 55.140 ;
        RECT 99.125 54.290 99.425 55.140 ;
        RECT 101.125 54.290 101.425 55.140 ;
        RECT 103.125 54.290 103.425 55.140 ;
        RECT 105.125 54.290 105.425 55.140 ;
        RECT 107.125 54.290 107.425 55.140 ;
        RECT 109.125 54.290 109.425 55.140 ;
        RECT 111.125 54.290 111.425 55.140 ;
        RECT 113.125 54.290 113.425 55.140 ;
        RECT 115.125 54.290 115.425 55.140 ;
        RECT 117.125 54.290 117.425 55.140 ;
        RECT 119.125 54.290 119.425 55.140 ;
        RECT 121.125 54.290 121.425 55.140 ;
        RECT 123.125 54.290 123.425 55.140 ;
        RECT 125.125 54.290 125.425 55.140 ;
        RECT 127.125 54.290 127.425 55.140 ;
        RECT 129.125 54.290 129.425 55.140 ;
        RECT 131.125 54.290 131.425 55.140 ;
        RECT 133.125 54.290 133.425 55.140 ;
        RECT 135.125 54.290 135.425 55.140 ;
        RECT 137.125 54.290 137.425 55.140 ;
        RECT 139.125 54.290 139.425 55.140 ;
        RECT 141.125 54.290 141.425 55.140 ;
        RECT 143.125 54.290 143.425 55.140 ;
        RECT 145.125 54.290 145.425 55.140 ;
        RECT 147.125 54.290 147.425 55.140 ;
        RECT 149.125 54.290 149.425 55.140 ;
        RECT 151.125 54.290 151.425 55.140 ;
        RECT 153.125 54.290 153.425 55.140 ;
        RECT 7.340 53.290 8.340 54.290 ;
        RECT 9.340 53.290 10.340 54.290 ;
        RECT 11.340 53.290 12.340 54.290 ;
        RECT 13.340 53.290 14.340 54.290 ;
        RECT 15.340 53.290 16.340 54.290 ;
        RECT 17.340 53.290 18.340 54.290 ;
        RECT 19.340 53.290 20.340 54.290 ;
        RECT 21.340 53.290 22.340 54.290 ;
        RECT 23.340 53.290 24.340 54.290 ;
        RECT 25.340 53.290 26.340 54.290 ;
        RECT 27.340 53.290 28.340 54.290 ;
        RECT 29.340 53.290 30.340 54.290 ;
        RECT 31.340 53.290 32.340 54.290 ;
        RECT 33.340 53.290 34.340 54.290 ;
        RECT 35.340 53.290 36.340 54.290 ;
        RECT 37.340 53.290 38.340 54.290 ;
        RECT 39.340 53.290 40.340 54.290 ;
        RECT 41.340 53.290 42.340 54.290 ;
        RECT 43.340 53.290 44.340 54.290 ;
        RECT 45.340 53.290 46.340 54.290 ;
        RECT 47.340 53.290 48.340 54.290 ;
        RECT 49.340 53.290 50.340 54.290 ;
        RECT 51.340 53.290 52.340 54.290 ;
        RECT 53.340 53.290 54.340 54.290 ;
        RECT 55.340 53.290 56.340 54.290 ;
        RECT 57.340 53.290 58.340 54.290 ;
        RECT 59.340 53.290 60.340 54.290 ;
        RECT 61.340 53.290 62.340 54.290 ;
        RECT 63.340 53.290 64.340 54.290 ;
        RECT 65.340 53.290 66.340 54.290 ;
        RECT 67.340 53.290 68.340 54.290 ;
        RECT 69.340 53.290 70.340 54.290 ;
        RECT 71.340 53.290 72.340 54.290 ;
        RECT 73.340 53.290 74.340 54.290 ;
        RECT 86.775 53.290 87.775 54.290 ;
        RECT 88.775 53.290 89.775 54.290 ;
        RECT 90.775 53.290 91.775 54.290 ;
        RECT 92.775 53.290 93.775 54.290 ;
        RECT 94.775 53.290 95.775 54.290 ;
        RECT 96.775 53.290 97.775 54.290 ;
        RECT 98.775 53.290 99.775 54.290 ;
        RECT 100.775 53.290 101.775 54.290 ;
        RECT 102.775 53.290 103.775 54.290 ;
        RECT 104.775 53.290 105.775 54.290 ;
        RECT 106.775 53.290 107.775 54.290 ;
        RECT 108.775 53.290 109.775 54.290 ;
        RECT 110.775 53.290 111.775 54.290 ;
        RECT 112.775 53.290 113.775 54.290 ;
        RECT 114.775 53.290 115.775 54.290 ;
        RECT 116.775 53.290 117.775 54.290 ;
        RECT 118.775 53.290 119.775 54.290 ;
        RECT 120.775 53.290 121.775 54.290 ;
        RECT 122.775 53.290 123.775 54.290 ;
        RECT 124.775 53.290 125.775 54.290 ;
        RECT 126.775 53.290 127.775 54.290 ;
        RECT 128.775 53.290 129.775 54.290 ;
        RECT 130.775 53.290 131.775 54.290 ;
        RECT 132.775 53.290 133.775 54.290 ;
        RECT 134.775 53.290 135.775 54.290 ;
        RECT 136.775 53.290 137.775 54.290 ;
        RECT 138.775 53.290 139.775 54.290 ;
        RECT 140.775 53.290 141.775 54.290 ;
        RECT 142.775 53.290 143.775 54.290 ;
        RECT 144.775 53.290 145.775 54.290 ;
        RECT 146.775 53.290 147.775 54.290 ;
        RECT 148.775 53.290 149.775 54.290 ;
        RECT 150.775 53.290 151.775 54.290 ;
        RECT 152.775 53.290 153.775 54.290 ;
        RECT 7.690 52.440 7.990 53.290 ;
        RECT 9.690 52.440 9.990 53.290 ;
        RECT 11.690 52.440 11.990 53.290 ;
        RECT 13.690 52.440 13.990 53.290 ;
        RECT 15.690 52.440 15.990 53.290 ;
        RECT 17.690 52.440 17.990 53.290 ;
        RECT 19.690 52.440 19.990 53.290 ;
        RECT 21.690 52.440 21.990 53.290 ;
        RECT 23.690 52.440 23.990 53.290 ;
        RECT 25.690 52.440 25.990 53.290 ;
        RECT 27.690 52.440 27.990 53.290 ;
        RECT 29.690 52.440 29.990 53.290 ;
        RECT 31.690 52.440 31.990 53.290 ;
        RECT 33.690 52.440 33.990 53.290 ;
        RECT 35.690 52.440 35.990 53.290 ;
        RECT 37.690 52.440 37.990 53.290 ;
        RECT 39.690 52.440 39.990 53.290 ;
        RECT 41.690 52.440 41.990 53.290 ;
        RECT 43.690 52.440 43.990 53.290 ;
        RECT 45.690 52.440 45.990 53.290 ;
        RECT 47.690 52.440 47.990 53.290 ;
        RECT 49.690 52.440 49.990 53.290 ;
        RECT 51.690 52.440 51.990 53.290 ;
        RECT 53.690 52.440 53.990 53.290 ;
        RECT 55.690 52.440 55.990 53.290 ;
        RECT 57.690 52.440 57.990 53.290 ;
        RECT 59.690 52.440 59.990 53.290 ;
        RECT 61.690 52.440 61.990 53.290 ;
        RECT 63.690 52.440 63.990 53.290 ;
        RECT 65.690 52.440 65.990 53.290 ;
        RECT 67.690 52.440 67.990 53.290 ;
        RECT 69.690 52.440 69.990 53.290 ;
        RECT 71.690 52.440 71.990 53.290 ;
        RECT 73.690 52.440 73.990 53.290 ;
        RECT 87.125 52.440 87.425 53.290 ;
        RECT 89.125 52.440 89.425 53.290 ;
        RECT 91.125 52.440 91.425 53.290 ;
        RECT 93.125 52.440 93.425 53.290 ;
        RECT 95.125 52.440 95.425 53.290 ;
        RECT 97.125 52.440 97.425 53.290 ;
        RECT 99.125 52.440 99.425 53.290 ;
        RECT 101.125 52.440 101.425 53.290 ;
        RECT 103.125 52.440 103.425 53.290 ;
        RECT 105.125 52.440 105.425 53.290 ;
        RECT 107.125 52.440 107.425 53.290 ;
        RECT 109.125 52.440 109.425 53.290 ;
        RECT 111.125 52.440 111.425 53.290 ;
        RECT 113.125 52.440 113.425 53.290 ;
        RECT 115.125 52.440 115.425 53.290 ;
        RECT 117.125 52.440 117.425 53.290 ;
        RECT 119.125 52.440 119.425 53.290 ;
        RECT 121.125 52.440 121.425 53.290 ;
        RECT 123.125 52.440 123.425 53.290 ;
        RECT 125.125 52.440 125.425 53.290 ;
        RECT 127.125 52.440 127.425 53.290 ;
        RECT 129.125 52.440 129.425 53.290 ;
        RECT 131.125 52.440 131.425 53.290 ;
        RECT 133.125 52.440 133.425 53.290 ;
        RECT 135.125 52.440 135.425 53.290 ;
        RECT 137.125 52.440 137.425 53.290 ;
        RECT 139.125 52.440 139.425 53.290 ;
        RECT 141.125 52.440 141.425 53.290 ;
        RECT 143.125 52.440 143.425 53.290 ;
        RECT 145.125 52.440 145.425 53.290 ;
        RECT 147.125 52.440 147.425 53.290 ;
        RECT 149.125 52.440 149.425 53.290 ;
        RECT 151.125 52.440 151.425 53.290 ;
        RECT 153.125 52.440 153.425 53.290 ;
        RECT 7.340 51.440 8.340 52.440 ;
        RECT 9.340 51.440 10.340 52.440 ;
        RECT 11.340 51.440 12.340 52.440 ;
        RECT 13.340 51.440 14.340 52.440 ;
        RECT 15.340 51.440 16.340 52.440 ;
        RECT 17.340 51.440 18.340 52.440 ;
        RECT 19.340 51.440 20.340 52.440 ;
        RECT 21.340 51.440 22.340 52.440 ;
        RECT 23.340 51.440 24.340 52.440 ;
        RECT 25.340 51.440 26.340 52.440 ;
        RECT 27.340 51.440 28.340 52.440 ;
        RECT 29.340 51.440 30.340 52.440 ;
        RECT 31.340 51.440 32.340 52.440 ;
        RECT 33.340 51.440 34.340 52.440 ;
        RECT 35.340 51.440 36.340 52.440 ;
        RECT 37.340 51.440 38.340 52.440 ;
        RECT 39.340 51.440 40.340 52.440 ;
        RECT 41.340 51.440 42.340 52.440 ;
        RECT 43.340 51.440 44.340 52.440 ;
        RECT 45.340 51.440 46.340 52.440 ;
        RECT 47.340 51.440 48.340 52.440 ;
        RECT 49.340 51.440 50.340 52.440 ;
        RECT 51.340 51.440 52.340 52.440 ;
        RECT 53.340 51.440 54.340 52.440 ;
        RECT 55.340 51.440 56.340 52.440 ;
        RECT 57.340 51.440 58.340 52.440 ;
        RECT 59.340 51.440 60.340 52.440 ;
        RECT 61.340 51.440 62.340 52.440 ;
        RECT 63.340 51.440 64.340 52.440 ;
        RECT 65.340 51.440 66.340 52.440 ;
        RECT 67.340 51.440 68.340 52.440 ;
        RECT 69.340 51.440 70.340 52.440 ;
        RECT 71.340 51.440 72.340 52.440 ;
        RECT 73.340 51.440 74.340 52.440 ;
        RECT 86.775 51.440 87.775 52.440 ;
        RECT 88.775 51.440 89.775 52.440 ;
        RECT 90.775 51.440 91.775 52.440 ;
        RECT 92.775 51.440 93.775 52.440 ;
        RECT 94.775 51.440 95.775 52.440 ;
        RECT 96.775 51.440 97.775 52.440 ;
        RECT 98.775 51.440 99.775 52.440 ;
        RECT 100.775 51.440 101.775 52.440 ;
        RECT 102.775 51.440 103.775 52.440 ;
        RECT 104.775 51.440 105.775 52.440 ;
        RECT 106.775 51.440 107.775 52.440 ;
        RECT 108.775 51.440 109.775 52.440 ;
        RECT 110.775 51.440 111.775 52.440 ;
        RECT 112.775 51.440 113.775 52.440 ;
        RECT 114.775 51.440 115.775 52.440 ;
        RECT 116.775 51.440 117.775 52.440 ;
        RECT 118.775 51.440 119.775 52.440 ;
        RECT 120.775 51.440 121.775 52.440 ;
        RECT 122.775 51.440 123.775 52.440 ;
        RECT 124.775 51.440 125.775 52.440 ;
        RECT 126.775 51.440 127.775 52.440 ;
        RECT 128.775 51.440 129.775 52.440 ;
        RECT 130.775 51.440 131.775 52.440 ;
        RECT 132.775 51.440 133.775 52.440 ;
        RECT 134.775 51.440 135.775 52.440 ;
        RECT 136.775 51.440 137.775 52.440 ;
        RECT 138.775 51.440 139.775 52.440 ;
        RECT 140.775 51.440 141.775 52.440 ;
        RECT 142.775 51.440 143.775 52.440 ;
        RECT 144.775 51.440 145.775 52.440 ;
        RECT 146.775 51.440 147.775 52.440 ;
        RECT 148.775 51.440 149.775 52.440 ;
        RECT 150.775 51.440 151.775 52.440 ;
        RECT 152.775 51.440 153.775 52.440 ;
        RECT 7.690 50.590 7.990 51.440 ;
        RECT 9.690 50.590 9.990 51.440 ;
        RECT 11.690 50.590 11.990 51.440 ;
        RECT 13.690 50.590 13.990 51.440 ;
        RECT 15.690 50.590 15.990 51.440 ;
        RECT 17.690 50.590 17.990 51.440 ;
        RECT 19.690 50.590 19.990 51.440 ;
        RECT 21.690 50.590 21.990 51.440 ;
        RECT 23.690 50.590 23.990 51.440 ;
        RECT 25.690 50.590 25.990 51.440 ;
        RECT 27.690 50.590 27.990 51.440 ;
        RECT 29.690 50.590 29.990 51.440 ;
        RECT 31.690 50.590 31.990 51.440 ;
        RECT 33.690 50.590 33.990 51.440 ;
        RECT 35.690 50.590 35.990 51.440 ;
        RECT 37.690 50.590 37.990 51.440 ;
        RECT 39.690 50.590 39.990 51.440 ;
        RECT 41.690 50.590 41.990 51.440 ;
        RECT 43.690 50.590 43.990 51.440 ;
        RECT 45.690 50.590 45.990 51.440 ;
        RECT 47.690 50.590 47.990 51.440 ;
        RECT 49.690 50.590 49.990 51.440 ;
        RECT 51.690 50.590 51.990 51.440 ;
        RECT 53.690 50.590 53.990 51.440 ;
        RECT 55.690 50.590 55.990 51.440 ;
        RECT 57.690 50.590 57.990 51.440 ;
        RECT 59.690 50.590 59.990 51.440 ;
        RECT 61.690 50.590 61.990 51.440 ;
        RECT 63.690 50.590 63.990 51.440 ;
        RECT 65.690 50.590 65.990 51.440 ;
        RECT 67.690 50.590 67.990 51.440 ;
        RECT 69.690 50.590 69.990 51.440 ;
        RECT 71.690 50.590 71.990 51.440 ;
        RECT 73.690 50.590 73.990 51.440 ;
        RECT 87.125 50.590 87.425 51.440 ;
        RECT 89.125 50.590 89.425 51.440 ;
        RECT 91.125 50.590 91.425 51.440 ;
        RECT 93.125 50.590 93.425 51.440 ;
        RECT 95.125 50.590 95.425 51.440 ;
        RECT 97.125 50.590 97.425 51.440 ;
        RECT 99.125 50.590 99.425 51.440 ;
        RECT 101.125 50.590 101.425 51.440 ;
        RECT 103.125 50.590 103.425 51.440 ;
        RECT 105.125 50.590 105.425 51.440 ;
        RECT 107.125 50.590 107.425 51.440 ;
        RECT 109.125 50.590 109.425 51.440 ;
        RECT 111.125 50.590 111.425 51.440 ;
        RECT 113.125 50.590 113.425 51.440 ;
        RECT 115.125 50.590 115.425 51.440 ;
        RECT 117.125 50.590 117.425 51.440 ;
        RECT 119.125 50.590 119.425 51.440 ;
        RECT 121.125 50.590 121.425 51.440 ;
        RECT 123.125 50.590 123.425 51.440 ;
        RECT 125.125 50.590 125.425 51.440 ;
        RECT 127.125 50.590 127.425 51.440 ;
        RECT 129.125 50.590 129.425 51.440 ;
        RECT 131.125 50.590 131.425 51.440 ;
        RECT 133.125 50.590 133.425 51.440 ;
        RECT 135.125 50.590 135.425 51.440 ;
        RECT 137.125 50.590 137.425 51.440 ;
        RECT 139.125 50.590 139.425 51.440 ;
        RECT 141.125 50.590 141.425 51.440 ;
        RECT 143.125 50.590 143.425 51.440 ;
        RECT 145.125 50.590 145.425 51.440 ;
        RECT 147.125 50.590 147.425 51.440 ;
        RECT 149.125 50.590 149.425 51.440 ;
        RECT 151.125 50.590 151.425 51.440 ;
        RECT 153.125 50.590 153.425 51.440 ;
        RECT 7.340 49.590 8.340 50.590 ;
        RECT 9.340 49.590 10.340 50.590 ;
        RECT 11.340 49.590 12.340 50.590 ;
        RECT 13.340 49.590 14.340 50.590 ;
        RECT 15.340 49.590 16.340 50.590 ;
        RECT 17.340 49.590 18.340 50.590 ;
        RECT 19.340 49.590 20.340 50.590 ;
        RECT 21.340 49.590 22.340 50.590 ;
        RECT 23.340 49.590 24.340 50.590 ;
        RECT 25.340 49.590 26.340 50.590 ;
        RECT 27.340 49.590 28.340 50.590 ;
        RECT 29.340 49.590 30.340 50.590 ;
        RECT 31.340 49.590 32.340 50.590 ;
        RECT 33.340 49.590 34.340 50.590 ;
        RECT 35.340 49.590 36.340 50.590 ;
        RECT 37.340 49.590 38.340 50.590 ;
        RECT 39.340 49.590 40.340 50.590 ;
        RECT 41.340 49.590 42.340 50.590 ;
        RECT 43.340 49.590 44.340 50.590 ;
        RECT 45.340 49.590 46.340 50.590 ;
        RECT 47.340 49.590 48.340 50.590 ;
        RECT 49.340 49.590 50.340 50.590 ;
        RECT 51.340 49.590 52.340 50.590 ;
        RECT 53.340 49.590 54.340 50.590 ;
        RECT 55.340 49.590 56.340 50.590 ;
        RECT 57.340 49.590 58.340 50.590 ;
        RECT 59.340 49.590 60.340 50.590 ;
        RECT 61.340 49.590 62.340 50.590 ;
        RECT 63.340 49.590 64.340 50.590 ;
        RECT 65.340 49.590 66.340 50.590 ;
        RECT 67.340 49.590 68.340 50.590 ;
        RECT 69.340 49.590 70.340 50.590 ;
        RECT 71.340 49.590 72.340 50.590 ;
        RECT 73.340 49.590 74.340 50.590 ;
        RECT 86.775 49.590 87.775 50.590 ;
        RECT 88.775 49.590 89.775 50.590 ;
        RECT 90.775 49.590 91.775 50.590 ;
        RECT 92.775 49.590 93.775 50.590 ;
        RECT 94.775 49.590 95.775 50.590 ;
        RECT 96.775 49.590 97.775 50.590 ;
        RECT 98.775 49.590 99.775 50.590 ;
        RECT 100.775 49.590 101.775 50.590 ;
        RECT 102.775 49.590 103.775 50.590 ;
        RECT 104.775 49.590 105.775 50.590 ;
        RECT 106.775 49.590 107.775 50.590 ;
        RECT 108.775 49.590 109.775 50.590 ;
        RECT 110.775 49.590 111.775 50.590 ;
        RECT 112.775 49.590 113.775 50.590 ;
        RECT 114.775 49.590 115.775 50.590 ;
        RECT 116.775 49.590 117.775 50.590 ;
        RECT 118.775 49.590 119.775 50.590 ;
        RECT 120.775 49.590 121.775 50.590 ;
        RECT 122.775 49.590 123.775 50.590 ;
        RECT 124.775 49.590 125.775 50.590 ;
        RECT 126.775 49.590 127.775 50.590 ;
        RECT 128.775 49.590 129.775 50.590 ;
        RECT 130.775 49.590 131.775 50.590 ;
        RECT 132.775 49.590 133.775 50.590 ;
        RECT 134.775 49.590 135.775 50.590 ;
        RECT 136.775 49.590 137.775 50.590 ;
        RECT 138.775 49.590 139.775 50.590 ;
        RECT 140.775 49.590 141.775 50.590 ;
        RECT 142.775 49.590 143.775 50.590 ;
        RECT 144.775 49.590 145.775 50.590 ;
        RECT 146.775 49.590 147.775 50.590 ;
        RECT 148.775 49.590 149.775 50.590 ;
        RECT 150.775 49.590 151.775 50.590 ;
        RECT 152.775 49.590 153.775 50.590 ;
        RECT 7.690 48.740 7.990 49.590 ;
        RECT 9.690 48.740 9.990 49.590 ;
        RECT 11.690 48.740 11.990 49.590 ;
        RECT 13.690 48.740 13.990 49.590 ;
        RECT 15.690 48.740 15.990 49.590 ;
        RECT 17.690 48.740 17.990 49.590 ;
        RECT 19.690 48.740 19.990 49.590 ;
        RECT 21.690 48.740 21.990 49.590 ;
        RECT 23.690 48.740 23.990 49.590 ;
        RECT 25.690 48.740 25.990 49.590 ;
        RECT 27.690 48.740 27.990 49.590 ;
        RECT 29.690 48.740 29.990 49.590 ;
        RECT 31.690 48.740 31.990 49.590 ;
        RECT 33.690 48.740 33.990 49.590 ;
        RECT 35.690 48.740 35.990 49.590 ;
        RECT 37.690 48.740 37.990 49.590 ;
        RECT 39.690 48.740 39.990 49.590 ;
        RECT 41.690 48.740 41.990 49.590 ;
        RECT 43.690 48.740 43.990 49.590 ;
        RECT 45.690 48.740 45.990 49.590 ;
        RECT 47.690 48.740 47.990 49.590 ;
        RECT 49.690 48.740 49.990 49.590 ;
        RECT 51.690 48.740 51.990 49.590 ;
        RECT 53.690 48.740 53.990 49.590 ;
        RECT 55.690 48.740 55.990 49.590 ;
        RECT 57.690 48.740 57.990 49.590 ;
        RECT 59.690 48.740 59.990 49.590 ;
        RECT 61.690 48.740 61.990 49.590 ;
        RECT 63.690 48.740 63.990 49.590 ;
        RECT 65.690 48.740 65.990 49.590 ;
        RECT 67.690 48.740 67.990 49.590 ;
        RECT 69.690 48.740 69.990 49.590 ;
        RECT 71.690 48.740 71.990 49.590 ;
        RECT 73.690 48.740 73.990 49.590 ;
        RECT 87.125 48.740 87.425 49.590 ;
        RECT 89.125 48.740 89.425 49.590 ;
        RECT 91.125 48.740 91.425 49.590 ;
        RECT 93.125 48.740 93.425 49.590 ;
        RECT 95.125 48.740 95.425 49.590 ;
        RECT 97.125 48.740 97.425 49.590 ;
        RECT 99.125 48.740 99.425 49.590 ;
        RECT 101.125 48.740 101.425 49.590 ;
        RECT 103.125 48.740 103.425 49.590 ;
        RECT 105.125 48.740 105.425 49.590 ;
        RECT 107.125 48.740 107.425 49.590 ;
        RECT 109.125 48.740 109.425 49.590 ;
        RECT 111.125 48.740 111.425 49.590 ;
        RECT 113.125 48.740 113.425 49.590 ;
        RECT 115.125 48.740 115.425 49.590 ;
        RECT 117.125 48.740 117.425 49.590 ;
        RECT 119.125 48.740 119.425 49.590 ;
        RECT 121.125 48.740 121.425 49.590 ;
        RECT 123.125 48.740 123.425 49.590 ;
        RECT 125.125 48.740 125.425 49.590 ;
        RECT 127.125 48.740 127.425 49.590 ;
        RECT 129.125 48.740 129.425 49.590 ;
        RECT 131.125 48.740 131.425 49.590 ;
        RECT 133.125 48.740 133.425 49.590 ;
        RECT 135.125 48.740 135.425 49.590 ;
        RECT 137.125 48.740 137.425 49.590 ;
        RECT 139.125 48.740 139.425 49.590 ;
        RECT 141.125 48.740 141.425 49.590 ;
        RECT 143.125 48.740 143.425 49.590 ;
        RECT 145.125 48.740 145.425 49.590 ;
        RECT 147.125 48.740 147.425 49.590 ;
        RECT 149.125 48.740 149.425 49.590 ;
        RECT 151.125 48.740 151.425 49.590 ;
        RECT 153.125 48.740 153.425 49.590 ;
        RECT 7.340 47.740 8.340 48.740 ;
        RECT 9.340 47.740 10.340 48.740 ;
        RECT 11.340 47.740 12.340 48.740 ;
        RECT 13.340 47.740 14.340 48.740 ;
        RECT 15.340 47.740 16.340 48.740 ;
        RECT 17.340 47.740 18.340 48.740 ;
        RECT 19.340 47.740 20.340 48.740 ;
        RECT 21.340 47.740 22.340 48.740 ;
        RECT 23.340 47.740 24.340 48.740 ;
        RECT 25.340 47.740 26.340 48.740 ;
        RECT 27.340 47.740 28.340 48.740 ;
        RECT 29.340 47.740 30.340 48.740 ;
        RECT 31.340 47.740 32.340 48.740 ;
        RECT 33.340 47.740 34.340 48.740 ;
        RECT 35.340 47.740 36.340 48.740 ;
        RECT 37.340 47.740 38.340 48.740 ;
        RECT 39.340 47.740 40.340 48.740 ;
        RECT 41.340 47.740 42.340 48.740 ;
        RECT 43.340 47.740 44.340 48.740 ;
        RECT 45.340 47.740 46.340 48.740 ;
        RECT 47.340 47.740 48.340 48.740 ;
        RECT 49.340 47.740 50.340 48.740 ;
        RECT 51.340 47.740 52.340 48.740 ;
        RECT 53.340 47.740 54.340 48.740 ;
        RECT 55.340 47.740 56.340 48.740 ;
        RECT 57.340 47.740 58.340 48.740 ;
        RECT 59.340 47.740 60.340 48.740 ;
        RECT 61.340 47.740 62.340 48.740 ;
        RECT 63.340 47.740 64.340 48.740 ;
        RECT 65.340 47.740 66.340 48.740 ;
        RECT 67.340 47.740 68.340 48.740 ;
        RECT 69.340 47.740 70.340 48.740 ;
        RECT 71.340 47.740 72.340 48.740 ;
        RECT 73.340 47.740 74.340 48.740 ;
        RECT 86.775 47.740 87.775 48.740 ;
        RECT 88.775 47.740 89.775 48.740 ;
        RECT 90.775 47.740 91.775 48.740 ;
        RECT 92.775 47.740 93.775 48.740 ;
        RECT 94.775 47.740 95.775 48.740 ;
        RECT 96.775 47.740 97.775 48.740 ;
        RECT 98.775 47.740 99.775 48.740 ;
        RECT 100.775 47.740 101.775 48.740 ;
        RECT 102.775 47.740 103.775 48.740 ;
        RECT 104.775 47.740 105.775 48.740 ;
        RECT 106.775 47.740 107.775 48.740 ;
        RECT 108.775 47.740 109.775 48.740 ;
        RECT 110.775 47.740 111.775 48.740 ;
        RECT 112.775 47.740 113.775 48.740 ;
        RECT 114.775 47.740 115.775 48.740 ;
        RECT 116.775 47.740 117.775 48.740 ;
        RECT 118.775 47.740 119.775 48.740 ;
        RECT 120.775 47.740 121.775 48.740 ;
        RECT 122.775 47.740 123.775 48.740 ;
        RECT 124.775 47.740 125.775 48.740 ;
        RECT 126.775 47.740 127.775 48.740 ;
        RECT 128.775 47.740 129.775 48.740 ;
        RECT 130.775 47.740 131.775 48.740 ;
        RECT 132.775 47.740 133.775 48.740 ;
        RECT 134.775 47.740 135.775 48.740 ;
        RECT 136.775 47.740 137.775 48.740 ;
        RECT 138.775 47.740 139.775 48.740 ;
        RECT 140.775 47.740 141.775 48.740 ;
        RECT 142.775 47.740 143.775 48.740 ;
        RECT 144.775 47.740 145.775 48.740 ;
        RECT 146.775 47.740 147.775 48.740 ;
        RECT 148.775 47.740 149.775 48.740 ;
        RECT 150.775 47.740 151.775 48.740 ;
        RECT 152.775 47.740 153.775 48.740 ;
        RECT 7.690 46.890 7.990 47.740 ;
        RECT 9.690 46.890 9.990 47.740 ;
        RECT 11.690 46.890 11.990 47.740 ;
        RECT 13.690 46.890 13.990 47.740 ;
        RECT 15.690 46.890 15.990 47.740 ;
        RECT 17.690 46.890 17.990 47.740 ;
        RECT 19.690 46.890 19.990 47.740 ;
        RECT 21.690 46.890 21.990 47.740 ;
        RECT 23.690 46.890 23.990 47.740 ;
        RECT 25.690 46.890 25.990 47.740 ;
        RECT 27.690 46.890 27.990 47.740 ;
        RECT 29.690 46.890 29.990 47.740 ;
        RECT 31.690 46.890 31.990 47.740 ;
        RECT 33.690 46.890 33.990 47.740 ;
        RECT 35.690 46.890 35.990 47.740 ;
        RECT 37.690 46.890 37.990 47.740 ;
        RECT 39.690 46.890 39.990 47.740 ;
        RECT 41.690 46.890 41.990 47.740 ;
        RECT 43.690 46.890 43.990 47.740 ;
        RECT 45.690 46.890 45.990 47.740 ;
        RECT 47.690 46.890 47.990 47.740 ;
        RECT 49.690 46.890 49.990 47.740 ;
        RECT 51.690 46.890 51.990 47.740 ;
        RECT 53.690 46.890 53.990 47.740 ;
        RECT 55.690 46.890 55.990 47.740 ;
        RECT 57.690 46.890 57.990 47.740 ;
        RECT 59.690 46.890 59.990 47.740 ;
        RECT 61.690 46.890 61.990 47.740 ;
        RECT 63.690 46.890 63.990 47.740 ;
        RECT 65.690 46.890 65.990 47.740 ;
        RECT 67.690 46.890 67.990 47.740 ;
        RECT 69.690 46.890 69.990 47.740 ;
        RECT 71.690 46.890 71.990 47.740 ;
        RECT 73.690 46.890 73.990 47.740 ;
        RECT 87.125 46.890 87.425 47.740 ;
        RECT 89.125 46.890 89.425 47.740 ;
        RECT 91.125 46.890 91.425 47.740 ;
        RECT 93.125 46.890 93.425 47.740 ;
        RECT 95.125 46.890 95.425 47.740 ;
        RECT 97.125 46.890 97.425 47.740 ;
        RECT 99.125 46.890 99.425 47.740 ;
        RECT 101.125 46.890 101.425 47.740 ;
        RECT 103.125 46.890 103.425 47.740 ;
        RECT 105.125 46.890 105.425 47.740 ;
        RECT 107.125 46.890 107.425 47.740 ;
        RECT 109.125 46.890 109.425 47.740 ;
        RECT 111.125 46.890 111.425 47.740 ;
        RECT 113.125 46.890 113.425 47.740 ;
        RECT 115.125 46.890 115.425 47.740 ;
        RECT 117.125 46.890 117.425 47.740 ;
        RECT 119.125 46.890 119.425 47.740 ;
        RECT 121.125 46.890 121.425 47.740 ;
        RECT 123.125 46.890 123.425 47.740 ;
        RECT 125.125 46.890 125.425 47.740 ;
        RECT 127.125 46.890 127.425 47.740 ;
        RECT 129.125 46.890 129.425 47.740 ;
        RECT 131.125 46.890 131.425 47.740 ;
        RECT 133.125 46.890 133.425 47.740 ;
        RECT 135.125 46.890 135.425 47.740 ;
        RECT 137.125 46.890 137.425 47.740 ;
        RECT 139.125 46.890 139.425 47.740 ;
        RECT 141.125 46.890 141.425 47.740 ;
        RECT 143.125 46.890 143.425 47.740 ;
        RECT 145.125 46.890 145.425 47.740 ;
        RECT 147.125 46.890 147.425 47.740 ;
        RECT 149.125 46.890 149.425 47.740 ;
        RECT 151.125 46.890 151.425 47.740 ;
        RECT 153.125 46.890 153.425 47.740 ;
        RECT 7.340 45.890 8.340 46.890 ;
        RECT 9.340 45.890 10.340 46.890 ;
        RECT 11.340 45.890 12.340 46.890 ;
        RECT 13.340 45.890 14.340 46.890 ;
        RECT 15.340 45.890 16.340 46.890 ;
        RECT 17.340 45.890 18.340 46.890 ;
        RECT 19.340 45.890 20.340 46.890 ;
        RECT 21.340 45.890 22.340 46.890 ;
        RECT 23.340 45.890 24.340 46.890 ;
        RECT 25.340 45.890 26.340 46.890 ;
        RECT 27.340 45.890 28.340 46.890 ;
        RECT 29.340 45.890 30.340 46.890 ;
        RECT 31.340 45.890 32.340 46.890 ;
        RECT 33.340 45.890 34.340 46.890 ;
        RECT 35.340 45.890 36.340 46.890 ;
        RECT 37.340 45.890 38.340 46.890 ;
        RECT 39.340 45.890 40.340 46.890 ;
        RECT 41.340 45.890 42.340 46.890 ;
        RECT 43.340 45.890 44.340 46.890 ;
        RECT 45.340 45.890 46.340 46.890 ;
        RECT 47.340 45.890 48.340 46.890 ;
        RECT 49.340 45.890 50.340 46.890 ;
        RECT 51.340 45.890 52.340 46.890 ;
        RECT 53.340 45.890 54.340 46.890 ;
        RECT 55.340 45.890 56.340 46.890 ;
        RECT 57.340 45.890 58.340 46.890 ;
        RECT 59.340 45.890 60.340 46.890 ;
        RECT 61.340 45.890 62.340 46.890 ;
        RECT 63.340 45.890 64.340 46.890 ;
        RECT 65.340 45.890 66.340 46.890 ;
        RECT 67.340 45.890 68.340 46.890 ;
        RECT 69.340 45.890 70.340 46.890 ;
        RECT 71.340 45.890 72.340 46.890 ;
        RECT 73.340 45.890 74.340 46.890 ;
        RECT 86.775 45.890 87.775 46.890 ;
        RECT 88.775 45.890 89.775 46.890 ;
        RECT 90.775 45.890 91.775 46.890 ;
        RECT 92.775 45.890 93.775 46.890 ;
        RECT 94.775 45.890 95.775 46.890 ;
        RECT 96.775 45.890 97.775 46.890 ;
        RECT 98.775 45.890 99.775 46.890 ;
        RECT 100.775 45.890 101.775 46.890 ;
        RECT 102.775 45.890 103.775 46.890 ;
        RECT 104.775 45.890 105.775 46.890 ;
        RECT 106.775 45.890 107.775 46.890 ;
        RECT 108.775 45.890 109.775 46.890 ;
        RECT 110.775 45.890 111.775 46.890 ;
        RECT 112.775 45.890 113.775 46.890 ;
        RECT 114.775 45.890 115.775 46.890 ;
        RECT 116.775 45.890 117.775 46.890 ;
        RECT 118.775 45.890 119.775 46.890 ;
        RECT 120.775 45.890 121.775 46.890 ;
        RECT 122.775 45.890 123.775 46.890 ;
        RECT 124.775 45.890 125.775 46.890 ;
        RECT 126.775 45.890 127.775 46.890 ;
        RECT 128.775 45.890 129.775 46.890 ;
        RECT 130.775 45.890 131.775 46.890 ;
        RECT 132.775 45.890 133.775 46.890 ;
        RECT 134.775 45.890 135.775 46.890 ;
        RECT 136.775 45.890 137.775 46.890 ;
        RECT 138.775 45.890 139.775 46.890 ;
        RECT 140.775 45.890 141.775 46.890 ;
        RECT 142.775 45.890 143.775 46.890 ;
        RECT 144.775 45.890 145.775 46.890 ;
        RECT 146.775 45.890 147.775 46.890 ;
        RECT 148.775 45.890 149.775 46.890 ;
        RECT 150.775 45.890 151.775 46.890 ;
        RECT 152.775 45.890 153.775 46.890 ;
        RECT 7.690 45.040 7.990 45.890 ;
        RECT 9.690 45.040 9.990 45.890 ;
        RECT 11.690 45.040 11.990 45.890 ;
        RECT 13.690 45.040 13.990 45.890 ;
        RECT 15.690 45.040 15.990 45.890 ;
        RECT 17.690 45.040 17.990 45.890 ;
        RECT 19.690 45.040 19.990 45.890 ;
        RECT 21.690 45.040 21.990 45.890 ;
        RECT 23.690 45.040 23.990 45.890 ;
        RECT 25.690 45.040 25.990 45.890 ;
        RECT 27.690 45.040 27.990 45.890 ;
        RECT 29.690 45.040 29.990 45.890 ;
        RECT 31.690 45.040 31.990 45.890 ;
        RECT 33.690 45.040 33.990 45.890 ;
        RECT 35.690 45.040 35.990 45.890 ;
        RECT 37.690 45.040 37.990 45.890 ;
        RECT 39.690 45.040 39.990 45.890 ;
        RECT 41.690 45.040 41.990 45.890 ;
        RECT 43.690 45.040 43.990 45.890 ;
        RECT 45.690 45.040 45.990 45.890 ;
        RECT 47.690 45.040 47.990 45.890 ;
        RECT 49.690 45.040 49.990 45.890 ;
        RECT 51.690 45.040 51.990 45.890 ;
        RECT 53.690 45.040 53.990 45.890 ;
        RECT 55.690 45.040 55.990 45.890 ;
        RECT 57.690 45.040 57.990 45.890 ;
        RECT 59.690 45.040 59.990 45.890 ;
        RECT 61.690 45.040 61.990 45.890 ;
        RECT 63.690 45.040 63.990 45.890 ;
        RECT 65.690 45.040 65.990 45.890 ;
        RECT 67.690 45.040 67.990 45.890 ;
        RECT 69.690 45.040 69.990 45.890 ;
        RECT 71.690 45.040 71.990 45.890 ;
        RECT 73.690 45.040 73.990 45.890 ;
        RECT 87.125 45.040 87.425 45.890 ;
        RECT 89.125 45.040 89.425 45.890 ;
        RECT 91.125 45.040 91.425 45.890 ;
        RECT 93.125 45.040 93.425 45.890 ;
        RECT 95.125 45.040 95.425 45.890 ;
        RECT 97.125 45.040 97.425 45.890 ;
        RECT 99.125 45.040 99.425 45.890 ;
        RECT 101.125 45.040 101.425 45.890 ;
        RECT 103.125 45.040 103.425 45.890 ;
        RECT 105.125 45.040 105.425 45.890 ;
        RECT 107.125 45.040 107.425 45.890 ;
        RECT 109.125 45.040 109.425 45.890 ;
        RECT 111.125 45.040 111.425 45.890 ;
        RECT 113.125 45.040 113.425 45.890 ;
        RECT 115.125 45.040 115.425 45.890 ;
        RECT 117.125 45.040 117.425 45.890 ;
        RECT 119.125 45.040 119.425 45.890 ;
        RECT 121.125 45.040 121.425 45.890 ;
        RECT 123.125 45.040 123.425 45.890 ;
        RECT 125.125 45.040 125.425 45.890 ;
        RECT 127.125 45.040 127.425 45.890 ;
        RECT 129.125 45.040 129.425 45.890 ;
        RECT 131.125 45.040 131.425 45.890 ;
        RECT 133.125 45.040 133.425 45.890 ;
        RECT 135.125 45.040 135.425 45.890 ;
        RECT 137.125 45.040 137.425 45.890 ;
        RECT 139.125 45.040 139.425 45.890 ;
        RECT 141.125 45.040 141.425 45.890 ;
        RECT 143.125 45.040 143.425 45.890 ;
        RECT 145.125 45.040 145.425 45.890 ;
        RECT 147.125 45.040 147.425 45.890 ;
        RECT 149.125 45.040 149.425 45.890 ;
        RECT 151.125 45.040 151.425 45.890 ;
        RECT 153.125 45.040 153.425 45.890 ;
        RECT 7.340 44.040 8.340 45.040 ;
        RECT 9.340 44.040 10.340 45.040 ;
        RECT 11.340 44.040 12.340 45.040 ;
        RECT 13.340 44.040 14.340 45.040 ;
        RECT 15.340 44.040 16.340 45.040 ;
        RECT 17.340 44.040 18.340 45.040 ;
        RECT 19.340 44.040 20.340 45.040 ;
        RECT 21.340 44.040 22.340 45.040 ;
        RECT 23.340 44.040 24.340 45.040 ;
        RECT 25.340 44.040 26.340 45.040 ;
        RECT 27.340 44.040 28.340 45.040 ;
        RECT 29.340 44.040 30.340 45.040 ;
        RECT 31.340 44.040 32.340 45.040 ;
        RECT 33.340 44.040 34.340 45.040 ;
        RECT 35.340 44.040 36.340 45.040 ;
        RECT 37.340 44.040 38.340 45.040 ;
        RECT 39.340 44.040 40.340 45.040 ;
        RECT 41.340 44.040 42.340 45.040 ;
        RECT 43.340 44.040 44.340 45.040 ;
        RECT 45.340 44.040 46.340 45.040 ;
        RECT 47.340 44.040 48.340 45.040 ;
        RECT 49.340 44.040 50.340 45.040 ;
        RECT 51.340 44.040 52.340 45.040 ;
        RECT 53.340 44.040 54.340 45.040 ;
        RECT 55.340 44.040 56.340 45.040 ;
        RECT 57.340 44.040 58.340 45.040 ;
        RECT 59.340 44.040 60.340 45.040 ;
        RECT 61.340 44.040 62.340 45.040 ;
        RECT 63.340 44.040 64.340 45.040 ;
        RECT 65.340 44.040 66.340 45.040 ;
        RECT 67.340 44.040 68.340 45.040 ;
        RECT 69.340 44.040 70.340 45.040 ;
        RECT 71.340 44.040 72.340 45.040 ;
        RECT 73.340 44.040 74.340 45.040 ;
        RECT 86.775 44.040 87.775 45.040 ;
        RECT 88.775 44.040 89.775 45.040 ;
        RECT 90.775 44.040 91.775 45.040 ;
        RECT 92.775 44.040 93.775 45.040 ;
        RECT 94.775 44.040 95.775 45.040 ;
        RECT 96.775 44.040 97.775 45.040 ;
        RECT 98.775 44.040 99.775 45.040 ;
        RECT 100.775 44.040 101.775 45.040 ;
        RECT 102.775 44.040 103.775 45.040 ;
        RECT 104.775 44.040 105.775 45.040 ;
        RECT 106.775 44.040 107.775 45.040 ;
        RECT 108.775 44.040 109.775 45.040 ;
        RECT 110.775 44.040 111.775 45.040 ;
        RECT 112.775 44.040 113.775 45.040 ;
        RECT 114.775 44.040 115.775 45.040 ;
        RECT 116.775 44.040 117.775 45.040 ;
        RECT 118.775 44.040 119.775 45.040 ;
        RECT 120.775 44.040 121.775 45.040 ;
        RECT 122.775 44.040 123.775 45.040 ;
        RECT 124.775 44.040 125.775 45.040 ;
        RECT 126.775 44.040 127.775 45.040 ;
        RECT 128.775 44.040 129.775 45.040 ;
        RECT 130.775 44.040 131.775 45.040 ;
        RECT 132.775 44.040 133.775 45.040 ;
        RECT 134.775 44.040 135.775 45.040 ;
        RECT 136.775 44.040 137.775 45.040 ;
        RECT 138.775 44.040 139.775 45.040 ;
        RECT 140.775 44.040 141.775 45.040 ;
        RECT 142.775 44.040 143.775 45.040 ;
        RECT 144.775 44.040 145.775 45.040 ;
        RECT 146.775 44.040 147.775 45.040 ;
        RECT 148.775 44.040 149.775 45.040 ;
        RECT 150.775 44.040 151.775 45.040 ;
        RECT 152.775 44.040 153.775 45.040 ;
        RECT 7.690 43.190 7.990 44.040 ;
        RECT 9.690 43.190 9.990 44.040 ;
        RECT 11.690 43.190 11.990 44.040 ;
        RECT 13.690 43.190 13.990 44.040 ;
        RECT 15.690 43.190 15.990 44.040 ;
        RECT 17.690 43.190 17.990 44.040 ;
        RECT 19.690 43.190 19.990 44.040 ;
        RECT 21.690 43.190 21.990 44.040 ;
        RECT 23.690 43.190 23.990 44.040 ;
        RECT 25.690 43.190 25.990 44.040 ;
        RECT 27.690 43.190 27.990 44.040 ;
        RECT 29.690 43.190 29.990 44.040 ;
        RECT 31.690 43.190 31.990 44.040 ;
        RECT 33.690 43.190 33.990 44.040 ;
        RECT 35.690 43.190 35.990 44.040 ;
        RECT 37.690 43.190 37.990 44.040 ;
        RECT 39.690 43.190 39.990 44.040 ;
        RECT 41.690 43.190 41.990 44.040 ;
        RECT 43.690 43.190 43.990 44.040 ;
        RECT 45.690 43.190 45.990 44.040 ;
        RECT 47.690 43.190 47.990 44.040 ;
        RECT 49.690 43.190 49.990 44.040 ;
        RECT 51.690 43.190 51.990 44.040 ;
        RECT 53.690 43.190 53.990 44.040 ;
        RECT 55.690 43.190 55.990 44.040 ;
        RECT 57.690 43.190 57.990 44.040 ;
        RECT 59.690 43.190 59.990 44.040 ;
        RECT 61.690 43.190 61.990 44.040 ;
        RECT 63.690 43.190 63.990 44.040 ;
        RECT 65.690 43.190 65.990 44.040 ;
        RECT 67.690 43.190 67.990 44.040 ;
        RECT 69.690 43.190 69.990 44.040 ;
        RECT 71.690 43.190 71.990 44.040 ;
        RECT 73.690 43.190 73.990 44.040 ;
        RECT 87.125 43.190 87.425 44.040 ;
        RECT 89.125 43.190 89.425 44.040 ;
        RECT 91.125 43.190 91.425 44.040 ;
        RECT 93.125 43.190 93.425 44.040 ;
        RECT 95.125 43.190 95.425 44.040 ;
        RECT 97.125 43.190 97.425 44.040 ;
        RECT 99.125 43.190 99.425 44.040 ;
        RECT 101.125 43.190 101.425 44.040 ;
        RECT 103.125 43.190 103.425 44.040 ;
        RECT 105.125 43.190 105.425 44.040 ;
        RECT 107.125 43.190 107.425 44.040 ;
        RECT 109.125 43.190 109.425 44.040 ;
        RECT 111.125 43.190 111.425 44.040 ;
        RECT 113.125 43.190 113.425 44.040 ;
        RECT 115.125 43.190 115.425 44.040 ;
        RECT 117.125 43.190 117.425 44.040 ;
        RECT 119.125 43.190 119.425 44.040 ;
        RECT 121.125 43.190 121.425 44.040 ;
        RECT 123.125 43.190 123.425 44.040 ;
        RECT 125.125 43.190 125.425 44.040 ;
        RECT 127.125 43.190 127.425 44.040 ;
        RECT 129.125 43.190 129.425 44.040 ;
        RECT 131.125 43.190 131.425 44.040 ;
        RECT 133.125 43.190 133.425 44.040 ;
        RECT 135.125 43.190 135.425 44.040 ;
        RECT 137.125 43.190 137.425 44.040 ;
        RECT 139.125 43.190 139.425 44.040 ;
        RECT 141.125 43.190 141.425 44.040 ;
        RECT 143.125 43.190 143.425 44.040 ;
        RECT 145.125 43.190 145.425 44.040 ;
        RECT 147.125 43.190 147.425 44.040 ;
        RECT 149.125 43.190 149.425 44.040 ;
        RECT 151.125 43.190 151.425 44.040 ;
        RECT 153.125 43.190 153.425 44.040 ;
        RECT 7.340 42.190 8.340 43.190 ;
        RECT 9.340 42.190 10.340 43.190 ;
        RECT 11.340 42.190 12.340 43.190 ;
        RECT 13.340 42.190 14.340 43.190 ;
        RECT 15.340 42.190 16.340 43.190 ;
        RECT 17.340 42.190 18.340 43.190 ;
        RECT 19.340 42.190 20.340 43.190 ;
        RECT 21.340 42.190 22.340 43.190 ;
        RECT 23.340 42.190 24.340 43.190 ;
        RECT 25.340 42.190 26.340 43.190 ;
        RECT 27.340 42.190 28.340 43.190 ;
        RECT 29.340 42.190 30.340 43.190 ;
        RECT 31.340 42.190 32.340 43.190 ;
        RECT 33.340 42.190 34.340 43.190 ;
        RECT 35.340 42.190 36.340 43.190 ;
        RECT 37.340 42.190 38.340 43.190 ;
        RECT 39.340 42.190 40.340 43.190 ;
        RECT 41.340 42.190 42.340 43.190 ;
        RECT 43.340 42.190 44.340 43.190 ;
        RECT 45.340 42.190 46.340 43.190 ;
        RECT 47.340 42.190 48.340 43.190 ;
        RECT 49.340 42.190 50.340 43.190 ;
        RECT 51.340 42.190 52.340 43.190 ;
        RECT 53.340 42.190 54.340 43.190 ;
        RECT 55.340 42.190 56.340 43.190 ;
        RECT 57.340 42.190 58.340 43.190 ;
        RECT 59.340 42.190 60.340 43.190 ;
        RECT 61.340 42.190 62.340 43.190 ;
        RECT 63.340 42.190 64.340 43.190 ;
        RECT 65.340 42.190 66.340 43.190 ;
        RECT 67.340 42.190 68.340 43.190 ;
        RECT 69.340 42.190 70.340 43.190 ;
        RECT 71.340 42.190 72.340 43.190 ;
        RECT 73.340 42.190 74.340 43.190 ;
        RECT 86.775 42.190 87.775 43.190 ;
        RECT 88.775 42.190 89.775 43.190 ;
        RECT 90.775 42.190 91.775 43.190 ;
        RECT 92.775 42.190 93.775 43.190 ;
        RECT 94.775 42.190 95.775 43.190 ;
        RECT 96.775 42.190 97.775 43.190 ;
        RECT 98.775 42.190 99.775 43.190 ;
        RECT 100.775 42.190 101.775 43.190 ;
        RECT 102.775 42.190 103.775 43.190 ;
        RECT 104.775 42.190 105.775 43.190 ;
        RECT 106.775 42.190 107.775 43.190 ;
        RECT 108.775 42.190 109.775 43.190 ;
        RECT 110.775 42.190 111.775 43.190 ;
        RECT 112.775 42.190 113.775 43.190 ;
        RECT 114.775 42.190 115.775 43.190 ;
        RECT 116.775 42.190 117.775 43.190 ;
        RECT 118.775 42.190 119.775 43.190 ;
        RECT 120.775 42.190 121.775 43.190 ;
        RECT 122.775 42.190 123.775 43.190 ;
        RECT 124.775 42.190 125.775 43.190 ;
        RECT 126.775 42.190 127.775 43.190 ;
        RECT 128.775 42.190 129.775 43.190 ;
        RECT 130.775 42.190 131.775 43.190 ;
        RECT 132.775 42.190 133.775 43.190 ;
        RECT 134.775 42.190 135.775 43.190 ;
        RECT 136.775 42.190 137.775 43.190 ;
        RECT 138.775 42.190 139.775 43.190 ;
        RECT 140.775 42.190 141.775 43.190 ;
        RECT 142.775 42.190 143.775 43.190 ;
        RECT 144.775 42.190 145.775 43.190 ;
        RECT 146.775 42.190 147.775 43.190 ;
        RECT 148.775 42.190 149.775 43.190 ;
        RECT 150.775 42.190 151.775 43.190 ;
        RECT 152.775 42.190 153.775 43.190 ;
        RECT 7.690 41.340 7.990 42.190 ;
        RECT 9.690 41.340 9.990 42.190 ;
        RECT 11.690 41.340 11.990 42.190 ;
        RECT 13.690 41.340 13.990 42.190 ;
        RECT 15.690 41.340 15.990 42.190 ;
        RECT 17.690 41.340 17.990 42.190 ;
        RECT 19.690 41.340 19.990 42.190 ;
        RECT 21.690 41.340 21.990 42.190 ;
        RECT 23.690 41.340 23.990 42.190 ;
        RECT 25.690 41.340 25.990 42.190 ;
        RECT 27.690 41.340 27.990 42.190 ;
        RECT 29.690 41.340 29.990 42.190 ;
        RECT 31.690 41.340 31.990 42.190 ;
        RECT 33.690 41.340 33.990 42.190 ;
        RECT 35.690 41.340 35.990 42.190 ;
        RECT 37.690 41.340 37.990 42.190 ;
        RECT 39.690 41.340 39.990 42.190 ;
        RECT 41.690 41.340 41.990 42.190 ;
        RECT 43.690 41.340 43.990 42.190 ;
        RECT 45.690 41.340 45.990 42.190 ;
        RECT 47.690 41.340 47.990 42.190 ;
        RECT 49.690 41.340 49.990 42.190 ;
        RECT 51.690 41.340 51.990 42.190 ;
        RECT 53.690 41.340 53.990 42.190 ;
        RECT 55.690 41.340 55.990 42.190 ;
        RECT 57.690 41.340 57.990 42.190 ;
        RECT 59.690 41.340 59.990 42.190 ;
        RECT 61.690 41.340 61.990 42.190 ;
        RECT 63.690 41.340 63.990 42.190 ;
        RECT 65.690 41.340 65.990 42.190 ;
        RECT 67.690 41.340 67.990 42.190 ;
        RECT 69.690 41.340 69.990 42.190 ;
        RECT 71.690 41.340 71.990 42.190 ;
        RECT 73.690 41.340 73.990 42.190 ;
        RECT 87.125 41.340 87.425 42.190 ;
        RECT 89.125 41.340 89.425 42.190 ;
        RECT 91.125 41.340 91.425 42.190 ;
        RECT 93.125 41.340 93.425 42.190 ;
        RECT 95.125 41.340 95.425 42.190 ;
        RECT 97.125 41.340 97.425 42.190 ;
        RECT 99.125 41.340 99.425 42.190 ;
        RECT 101.125 41.340 101.425 42.190 ;
        RECT 103.125 41.340 103.425 42.190 ;
        RECT 105.125 41.340 105.425 42.190 ;
        RECT 107.125 41.340 107.425 42.190 ;
        RECT 109.125 41.340 109.425 42.190 ;
        RECT 111.125 41.340 111.425 42.190 ;
        RECT 113.125 41.340 113.425 42.190 ;
        RECT 115.125 41.340 115.425 42.190 ;
        RECT 117.125 41.340 117.425 42.190 ;
        RECT 119.125 41.340 119.425 42.190 ;
        RECT 121.125 41.340 121.425 42.190 ;
        RECT 123.125 41.340 123.425 42.190 ;
        RECT 125.125 41.340 125.425 42.190 ;
        RECT 127.125 41.340 127.425 42.190 ;
        RECT 129.125 41.340 129.425 42.190 ;
        RECT 131.125 41.340 131.425 42.190 ;
        RECT 133.125 41.340 133.425 42.190 ;
        RECT 135.125 41.340 135.425 42.190 ;
        RECT 137.125 41.340 137.425 42.190 ;
        RECT 139.125 41.340 139.425 42.190 ;
        RECT 141.125 41.340 141.425 42.190 ;
        RECT 143.125 41.340 143.425 42.190 ;
        RECT 145.125 41.340 145.425 42.190 ;
        RECT 147.125 41.340 147.425 42.190 ;
        RECT 149.125 41.340 149.425 42.190 ;
        RECT 151.125 41.340 151.425 42.190 ;
        RECT 153.125 41.340 153.425 42.190 ;
        RECT 7.340 40.340 8.340 41.340 ;
        RECT 9.340 40.340 10.340 41.340 ;
        RECT 11.340 40.340 12.340 41.340 ;
        RECT 13.340 40.340 14.340 41.340 ;
        RECT 15.340 40.340 16.340 41.340 ;
        RECT 17.340 40.340 18.340 41.340 ;
        RECT 19.340 40.340 20.340 41.340 ;
        RECT 21.340 40.340 22.340 41.340 ;
        RECT 23.340 40.340 24.340 41.340 ;
        RECT 25.340 40.340 26.340 41.340 ;
        RECT 27.340 40.340 28.340 41.340 ;
        RECT 29.340 40.340 30.340 41.340 ;
        RECT 31.340 40.340 32.340 41.340 ;
        RECT 33.340 40.340 34.340 41.340 ;
        RECT 35.340 40.340 36.340 41.340 ;
        RECT 37.340 40.340 38.340 41.340 ;
        RECT 39.340 40.340 40.340 41.340 ;
        RECT 41.340 40.340 42.340 41.340 ;
        RECT 43.340 40.340 44.340 41.340 ;
        RECT 45.340 40.340 46.340 41.340 ;
        RECT 47.340 40.340 48.340 41.340 ;
        RECT 49.340 40.340 50.340 41.340 ;
        RECT 51.340 40.340 52.340 41.340 ;
        RECT 53.340 40.340 54.340 41.340 ;
        RECT 55.340 40.340 56.340 41.340 ;
        RECT 57.340 40.340 58.340 41.340 ;
        RECT 59.340 40.340 60.340 41.340 ;
        RECT 61.340 40.340 62.340 41.340 ;
        RECT 63.340 40.340 64.340 41.340 ;
        RECT 65.340 40.340 66.340 41.340 ;
        RECT 67.340 40.340 68.340 41.340 ;
        RECT 69.340 40.340 70.340 41.340 ;
        RECT 71.340 40.340 72.340 41.340 ;
        RECT 73.340 40.340 74.340 41.340 ;
        RECT 86.775 40.340 87.775 41.340 ;
        RECT 88.775 40.340 89.775 41.340 ;
        RECT 90.775 40.340 91.775 41.340 ;
        RECT 92.775 40.340 93.775 41.340 ;
        RECT 94.775 40.340 95.775 41.340 ;
        RECT 96.775 40.340 97.775 41.340 ;
        RECT 98.775 40.340 99.775 41.340 ;
        RECT 100.775 40.340 101.775 41.340 ;
        RECT 102.775 40.340 103.775 41.340 ;
        RECT 104.775 40.340 105.775 41.340 ;
        RECT 106.775 40.340 107.775 41.340 ;
        RECT 108.775 40.340 109.775 41.340 ;
        RECT 110.775 40.340 111.775 41.340 ;
        RECT 112.775 40.340 113.775 41.340 ;
        RECT 114.775 40.340 115.775 41.340 ;
        RECT 116.775 40.340 117.775 41.340 ;
        RECT 118.775 40.340 119.775 41.340 ;
        RECT 120.775 40.340 121.775 41.340 ;
        RECT 122.775 40.340 123.775 41.340 ;
        RECT 124.775 40.340 125.775 41.340 ;
        RECT 126.775 40.340 127.775 41.340 ;
        RECT 128.775 40.340 129.775 41.340 ;
        RECT 130.775 40.340 131.775 41.340 ;
        RECT 132.775 40.340 133.775 41.340 ;
        RECT 134.775 40.340 135.775 41.340 ;
        RECT 136.775 40.340 137.775 41.340 ;
        RECT 138.775 40.340 139.775 41.340 ;
        RECT 140.775 40.340 141.775 41.340 ;
        RECT 142.775 40.340 143.775 41.340 ;
        RECT 144.775 40.340 145.775 41.340 ;
        RECT 146.775 40.340 147.775 41.340 ;
        RECT 148.775 40.340 149.775 41.340 ;
        RECT 150.775 40.340 151.775 41.340 ;
        RECT 152.775 40.340 153.775 41.340 ;
        RECT 7.690 39.490 7.990 40.340 ;
        RECT 9.690 39.490 9.990 40.340 ;
        RECT 11.690 39.490 11.990 40.340 ;
        RECT 13.690 39.490 13.990 40.340 ;
        RECT 15.690 39.490 15.990 40.340 ;
        RECT 17.690 39.490 17.990 40.340 ;
        RECT 19.690 39.490 19.990 40.340 ;
        RECT 21.690 39.490 21.990 40.340 ;
        RECT 23.690 39.490 23.990 40.340 ;
        RECT 25.690 39.490 25.990 40.340 ;
        RECT 27.690 39.490 27.990 40.340 ;
        RECT 29.690 39.490 29.990 40.340 ;
        RECT 31.690 39.490 31.990 40.340 ;
        RECT 33.690 39.490 33.990 40.340 ;
        RECT 35.690 39.490 35.990 40.340 ;
        RECT 37.690 39.490 37.990 40.340 ;
        RECT 39.690 39.490 39.990 40.340 ;
        RECT 41.690 39.490 41.990 40.340 ;
        RECT 43.690 39.490 43.990 40.340 ;
        RECT 45.690 39.490 45.990 40.340 ;
        RECT 47.690 39.490 47.990 40.340 ;
        RECT 49.690 39.490 49.990 40.340 ;
        RECT 51.690 39.490 51.990 40.340 ;
        RECT 53.690 39.490 53.990 40.340 ;
        RECT 55.690 39.490 55.990 40.340 ;
        RECT 57.690 39.490 57.990 40.340 ;
        RECT 59.690 39.490 59.990 40.340 ;
        RECT 61.690 39.490 61.990 40.340 ;
        RECT 63.690 39.490 63.990 40.340 ;
        RECT 65.690 39.490 65.990 40.340 ;
        RECT 67.690 39.490 67.990 40.340 ;
        RECT 69.690 39.490 69.990 40.340 ;
        RECT 71.690 39.490 71.990 40.340 ;
        RECT 73.690 39.490 73.990 40.340 ;
        RECT 87.125 39.490 87.425 40.340 ;
        RECT 89.125 39.490 89.425 40.340 ;
        RECT 91.125 39.490 91.425 40.340 ;
        RECT 93.125 39.490 93.425 40.340 ;
        RECT 95.125 39.490 95.425 40.340 ;
        RECT 97.125 39.490 97.425 40.340 ;
        RECT 99.125 39.490 99.425 40.340 ;
        RECT 101.125 39.490 101.425 40.340 ;
        RECT 103.125 39.490 103.425 40.340 ;
        RECT 105.125 39.490 105.425 40.340 ;
        RECT 107.125 39.490 107.425 40.340 ;
        RECT 109.125 39.490 109.425 40.340 ;
        RECT 111.125 39.490 111.425 40.340 ;
        RECT 113.125 39.490 113.425 40.340 ;
        RECT 115.125 39.490 115.425 40.340 ;
        RECT 117.125 39.490 117.425 40.340 ;
        RECT 119.125 39.490 119.425 40.340 ;
        RECT 121.125 39.490 121.425 40.340 ;
        RECT 123.125 39.490 123.425 40.340 ;
        RECT 125.125 39.490 125.425 40.340 ;
        RECT 127.125 39.490 127.425 40.340 ;
        RECT 129.125 39.490 129.425 40.340 ;
        RECT 131.125 39.490 131.425 40.340 ;
        RECT 133.125 39.490 133.425 40.340 ;
        RECT 135.125 39.490 135.425 40.340 ;
        RECT 137.125 39.490 137.425 40.340 ;
        RECT 139.125 39.490 139.425 40.340 ;
        RECT 141.125 39.490 141.425 40.340 ;
        RECT 143.125 39.490 143.425 40.340 ;
        RECT 145.125 39.490 145.425 40.340 ;
        RECT 147.125 39.490 147.425 40.340 ;
        RECT 149.125 39.490 149.425 40.340 ;
        RECT 151.125 39.490 151.425 40.340 ;
        RECT 153.125 39.490 153.425 40.340 ;
        RECT 7.340 38.490 8.340 39.490 ;
        RECT 9.340 38.490 10.340 39.490 ;
        RECT 11.340 38.490 12.340 39.490 ;
        RECT 13.340 38.490 14.340 39.490 ;
        RECT 15.340 38.490 16.340 39.490 ;
        RECT 17.340 38.490 18.340 39.490 ;
        RECT 19.340 38.490 20.340 39.490 ;
        RECT 21.340 38.490 22.340 39.490 ;
        RECT 23.340 38.490 24.340 39.490 ;
        RECT 25.340 38.490 26.340 39.490 ;
        RECT 27.340 38.490 28.340 39.490 ;
        RECT 29.340 38.490 30.340 39.490 ;
        RECT 31.340 38.490 32.340 39.490 ;
        RECT 33.340 38.490 34.340 39.490 ;
        RECT 35.340 38.490 36.340 39.490 ;
        RECT 37.340 38.490 38.340 39.490 ;
        RECT 39.340 38.490 40.340 39.490 ;
        RECT 41.340 38.490 42.340 39.490 ;
        RECT 43.340 38.490 44.340 39.490 ;
        RECT 45.340 38.490 46.340 39.490 ;
        RECT 47.340 38.490 48.340 39.490 ;
        RECT 49.340 38.490 50.340 39.490 ;
        RECT 51.340 38.490 52.340 39.490 ;
        RECT 53.340 38.490 54.340 39.490 ;
        RECT 55.340 38.490 56.340 39.490 ;
        RECT 57.340 38.490 58.340 39.490 ;
        RECT 59.340 38.490 60.340 39.490 ;
        RECT 61.340 38.490 62.340 39.490 ;
        RECT 63.340 38.490 64.340 39.490 ;
        RECT 65.340 38.490 66.340 39.490 ;
        RECT 67.340 38.490 68.340 39.490 ;
        RECT 69.340 38.490 70.340 39.490 ;
        RECT 71.340 38.490 72.340 39.490 ;
        RECT 73.340 38.490 74.340 39.490 ;
        RECT 86.775 38.490 87.775 39.490 ;
        RECT 88.775 38.490 89.775 39.490 ;
        RECT 90.775 38.490 91.775 39.490 ;
        RECT 92.775 38.490 93.775 39.490 ;
        RECT 94.775 38.490 95.775 39.490 ;
        RECT 96.775 38.490 97.775 39.490 ;
        RECT 98.775 38.490 99.775 39.490 ;
        RECT 100.775 38.490 101.775 39.490 ;
        RECT 102.775 38.490 103.775 39.490 ;
        RECT 104.775 38.490 105.775 39.490 ;
        RECT 106.775 38.490 107.775 39.490 ;
        RECT 108.775 38.490 109.775 39.490 ;
        RECT 110.775 38.490 111.775 39.490 ;
        RECT 112.775 38.490 113.775 39.490 ;
        RECT 114.775 38.490 115.775 39.490 ;
        RECT 116.775 38.490 117.775 39.490 ;
        RECT 118.775 38.490 119.775 39.490 ;
        RECT 120.775 38.490 121.775 39.490 ;
        RECT 122.775 38.490 123.775 39.490 ;
        RECT 124.775 38.490 125.775 39.490 ;
        RECT 126.775 38.490 127.775 39.490 ;
        RECT 128.775 38.490 129.775 39.490 ;
        RECT 130.775 38.490 131.775 39.490 ;
        RECT 132.775 38.490 133.775 39.490 ;
        RECT 134.775 38.490 135.775 39.490 ;
        RECT 136.775 38.490 137.775 39.490 ;
        RECT 138.775 38.490 139.775 39.490 ;
        RECT 140.775 38.490 141.775 39.490 ;
        RECT 142.775 38.490 143.775 39.490 ;
        RECT 144.775 38.490 145.775 39.490 ;
        RECT 146.775 38.490 147.775 39.490 ;
        RECT 148.775 38.490 149.775 39.490 ;
        RECT 150.775 38.490 151.775 39.490 ;
        RECT 152.775 38.490 153.775 39.490 ;
        RECT 7.690 37.640 7.990 38.490 ;
        RECT 9.690 37.640 9.990 38.490 ;
        RECT 11.690 37.640 11.990 38.490 ;
        RECT 13.690 37.640 13.990 38.490 ;
        RECT 15.690 37.640 15.990 38.490 ;
        RECT 17.690 37.640 17.990 38.490 ;
        RECT 19.690 37.640 19.990 38.490 ;
        RECT 21.690 37.640 21.990 38.490 ;
        RECT 23.690 37.640 23.990 38.490 ;
        RECT 25.690 37.640 25.990 38.490 ;
        RECT 27.690 37.640 27.990 38.490 ;
        RECT 29.690 37.640 29.990 38.490 ;
        RECT 31.690 37.640 31.990 38.490 ;
        RECT 33.690 37.640 33.990 38.490 ;
        RECT 35.690 37.640 35.990 38.490 ;
        RECT 37.690 37.640 37.990 38.490 ;
        RECT 39.690 37.640 39.990 38.490 ;
        RECT 41.690 37.640 41.990 38.490 ;
        RECT 43.690 37.640 43.990 38.490 ;
        RECT 45.690 37.640 45.990 38.490 ;
        RECT 47.690 37.640 47.990 38.490 ;
        RECT 49.690 37.640 49.990 38.490 ;
        RECT 51.690 37.640 51.990 38.490 ;
        RECT 53.690 37.640 53.990 38.490 ;
        RECT 55.690 37.640 55.990 38.490 ;
        RECT 57.690 37.640 57.990 38.490 ;
        RECT 59.690 37.640 59.990 38.490 ;
        RECT 61.690 37.640 61.990 38.490 ;
        RECT 63.690 37.640 63.990 38.490 ;
        RECT 65.690 37.640 65.990 38.490 ;
        RECT 67.690 37.640 67.990 38.490 ;
        RECT 69.690 37.640 69.990 38.490 ;
        RECT 71.690 37.640 71.990 38.490 ;
        RECT 73.690 37.640 73.990 38.490 ;
        RECT 87.125 37.640 87.425 38.490 ;
        RECT 89.125 37.640 89.425 38.490 ;
        RECT 91.125 37.640 91.425 38.490 ;
        RECT 93.125 37.640 93.425 38.490 ;
        RECT 95.125 37.640 95.425 38.490 ;
        RECT 97.125 37.640 97.425 38.490 ;
        RECT 99.125 37.640 99.425 38.490 ;
        RECT 101.125 37.640 101.425 38.490 ;
        RECT 103.125 37.640 103.425 38.490 ;
        RECT 105.125 37.640 105.425 38.490 ;
        RECT 107.125 37.640 107.425 38.490 ;
        RECT 109.125 37.640 109.425 38.490 ;
        RECT 111.125 37.640 111.425 38.490 ;
        RECT 113.125 37.640 113.425 38.490 ;
        RECT 115.125 37.640 115.425 38.490 ;
        RECT 117.125 37.640 117.425 38.490 ;
        RECT 119.125 37.640 119.425 38.490 ;
        RECT 121.125 37.640 121.425 38.490 ;
        RECT 123.125 37.640 123.425 38.490 ;
        RECT 125.125 37.640 125.425 38.490 ;
        RECT 127.125 37.640 127.425 38.490 ;
        RECT 129.125 37.640 129.425 38.490 ;
        RECT 131.125 37.640 131.425 38.490 ;
        RECT 133.125 37.640 133.425 38.490 ;
        RECT 135.125 37.640 135.425 38.490 ;
        RECT 137.125 37.640 137.425 38.490 ;
        RECT 139.125 37.640 139.425 38.490 ;
        RECT 141.125 37.640 141.425 38.490 ;
        RECT 143.125 37.640 143.425 38.490 ;
        RECT 145.125 37.640 145.425 38.490 ;
        RECT 147.125 37.640 147.425 38.490 ;
        RECT 149.125 37.640 149.425 38.490 ;
        RECT 151.125 37.640 151.425 38.490 ;
        RECT 153.125 37.640 153.425 38.490 ;
        RECT 7.340 36.640 8.340 37.640 ;
        RECT 9.340 36.640 10.340 37.640 ;
        RECT 11.340 36.640 12.340 37.640 ;
        RECT 13.340 36.640 14.340 37.640 ;
        RECT 15.340 36.640 16.340 37.640 ;
        RECT 17.340 36.640 18.340 37.640 ;
        RECT 19.340 36.640 20.340 37.640 ;
        RECT 21.340 36.640 22.340 37.640 ;
        RECT 23.340 36.640 24.340 37.640 ;
        RECT 25.340 36.640 26.340 37.640 ;
        RECT 27.340 36.640 28.340 37.640 ;
        RECT 29.340 36.640 30.340 37.640 ;
        RECT 31.340 36.640 32.340 37.640 ;
        RECT 33.340 36.640 34.340 37.640 ;
        RECT 35.340 36.640 36.340 37.640 ;
        RECT 37.340 36.640 38.340 37.640 ;
        RECT 39.340 36.640 40.340 37.640 ;
        RECT 41.340 36.640 42.340 37.640 ;
        RECT 43.340 36.640 44.340 37.640 ;
        RECT 45.340 36.640 46.340 37.640 ;
        RECT 47.340 36.640 48.340 37.640 ;
        RECT 49.340 36.640 50.340 37.640 ;
        RECT 51.340 36.640 52.340 37.640 ;
        RECT 53.340 36.640 54.340 37.640 ;
        RECT 55.340 36.640 56.340 37.640 ;
        RECT 57.340 36.640 58.340 37.640 ;
        RECT 59.340 36.640 60.340 37.640 ;
        RECT 61.340 36.640 62.340 37.640 ;
        RECT 63.340 36.640 64.340 37.640 ;
        RECT 65.340 36.640 66.340 37.640 ;
        RECT 67.340 36.640 68.340 37.640 ;
        RECT 69.340 36.640 70.340 37.640 ;
        RECT 71.340 36.640 72.340 37.640 ;
        RECT 73.340 36.640 74.340 37.640 ;
        RECT 86.775 36.640 87.775 37.640 ;
        RECT 88.775 36.640 89.775 37.640 ;
        RECT 90.775 36.640 91.775 37.640 ;
        RECT 92.775 36.640 93.775 37.640 ;
        RECT 94.775 36.640 95.775 37.640 ;
        RECT 96.775 36.640 97.775 37.640 ;
        RECT 98.775 36.640 99.775 37.640 ;
        RECT 100.775 36.640 101.775 37.640 ;
        RECT 102.775 36.640 103.775 37.640 ;
        RECT 104.775 36.640 105.775 37.640 ;
        RECT 106.775 36.640 107.775 37.640 ;
        RECT 108.775 36.640 109.775 37.640 ;
        RECT 110.775 36.640 111.775 37.640 ;
        RECT 112.775 36.640 113.775 37.640 ;
        RECT 114.775 36.640 115.775 37.640 ;
        RECT 116.775 36.640 117.775 37.640 ;
        RECT 118.775 36.640 119.775 37.640 ;
        RECT 120.775 36.640 121.775 37.640 ;
        RECT 122.775 36.640 123.775 37.640 ;
        RECT 124.775 36.640 125.775 37.640 ;
        RECT 126.775 36.640 127.775 37.640 ;
        RECT 128.775 36.640 129.775 37.640 ;
        RECT 130.775 36.640 131.775 37.640 ;
        RECT 132.775 36.640 133.775 37.640 ;
        RECT 134.775 36.640 135.775 37.640 ;
        RECT 136.775 36.640 137.775 37.640 ;
        RECT 138.775 36.640 139.775 37.640 ;
        RECT 140.775 36.640 141.775 37.640 ;
        RECT 142.775 36.640 143.775 37.640 ;
        RECT 144.775 36.640 145.775 37.640 ;
        RECT 146.775 36.640 147.775 37.640 ;
        RECT 148.775 36.640 149.775 37.640 ;
        RECT 150.775 36.640 151.775 37.640 ;
        RECT 152.775 36.640 153.775 37.640 ;
        RECT 7.690 35.790 7.990 36.640 ;
        RECT 9.690 35.790 9.990 36.640 ;
        RECT 11.690 35.790 11.990 36.640 ;
        RECT 13.690 35.790 13.990 36.640 ;
        RECT 15.690 35.790 15.990 36.640 ;
        RECT 17.690 35.790 17.990 36.640 ;
        RECT 19.690 35.790 19.990 36.640 ;
        RECT 21.690 35.790 21.990 36.640 ;
        RECT 23.690 35.790 23.990 36.640 ;
        RECT 25.690 35.790 25.990 36.640 ;
        RECT 27.690 35.790 27.990 36.640 ;
        RECT 29.690 35.790 29.990 36.640 ;
        RECT 31.690 35.790 31.990 36.640 ;
        RECT 33.690 35.790 33.990 36.640 ;
        RECT 35.690 35.790 35.990 36.640 ;
        RECT 37.690 35.790 37.990 36.640 ;
        RECT 39.690 35.790 39.990 36.640 ;
        RECT 41.690 35.790 41.990 36.640 ;
        RECT 43.690 35.790 43.990 36.640 ;
        RECT 45.690 35.790 45.990 36.640 ;
        RECT 47.690 35.790 47.990 36.640 ;
        RECT 49.690 35.790 49.990 36.640 ;
        RECT 51.690 35.790 51.990 36.640 ;
        RECT 53.690 35.790 53.990 36.640 ;
        RECT 55.690 35.790 55.990 36.640 ;
        RECT 57.690 35.790 57.990 36.640 ;
        RECT 59.690 35.790 59.990 36.640 ;
        RECT 61.690 35.790 61.990 36.640 ;
        RECT 63.690 35.790 63.990 36.640 ;
        RECT 65.690 35.790 65.990 36.640 ;
        RECT 67.690 35.790 67.990 36.640 ;
        RECT 69.690 35.790 69.990 36.640 ;
        RECT 71.690 35.790 71.990 36.640 ;
        RECT 73.690 35.790 73.990 36.640 ;
        RECT 87.125 35.790 87.425 36.640 ;
        RECT 89.125 35.790 89.425 36.640 ;
        RECT 91.125 35.790 91.425 36.640 ;
        RECT 93.125 35.790 93.425 36.640 ;
        RECT 95.125 35.790 95.425 36.640 ;
        RECT 97.125 35.790 97.425 36.640 ;
        RECT 99.125 35.790 99.425 36.640 ;
        RECT 101.125 35.790 101.425 36.640 ;
        RECT 103.125 35.790 103.425 36.640 ;
        RECT 105.125 35.790 105.425 36.640 ;
        RECT 107.125 35.790 107.425 36.640 ;
        RECT 109.125 35.790 109.425 36.640 ;
        RECT 111.125 35.790 111.425 36.640 ;
        RECT 113.125 35.790 113.425 36.640 ;
        RECT 115.125 35.790 115.425 36.640 ;
        RECT 117.125 35.790 117.425 36.640 ;
        RECT 119.125 35.790 119.425 36.640 ;
        RECT 121.125 35.790 121.425 36.640 ;
        RECT 123.125 35.790 123.425 36.640 ;
        RECT 125.125 35.790 125.425 36.640 ;
        RECT 127.125 35.790 127.425 36.640 ;
        RECT 129.125 35.790 129.425 36.640 ;
        RECT 131.125 35.790 131.425 36.640 ;
        RECT 133.125 35.790 133.425 36.640 ;
        RECT 135.125 35.790 135.425 36.640 ;
        RECT 137.125 35.790 137.425 36.640 ;
        RECT 139.125 35.790 139.425 36.640 ;
        RECT 141.125 35.790 141.425 36.640 ;
        RECT 143.125 35.790 143.425 36.640 ;
        RECT 145.125 35.790 145.425 36.640 ;
        RECT 147.125 35.790 147.425 36.640 ;
        RECT 149.125 35.790 149.425 36.640 ;
        RECT 151.125 35.790 151.425 36.640 ;
        RECT 153.125 35.790 153.425 36.640 ;
        RECT 7.340 34.790 8.340 35.790 ;
        RECT 9.340 34.790 10.340 35.790 ;
        RECT 11.340 34.790 12.340 35.790 ;
        RECT 13.340 34.790 14.340 35.790 ;
        RECT 15.340 34.790 16.340 35.790 ;
        RECT 17.340 34.790 18.340 35.790 ;
        RECT 19.340 34.790 20.340 35.790 ;
        RECT 21.340 34.790 22.340 35.790 ;
        RECT 23.340 34.790 24.340 35.790 ;
        RECT 25.340 34.790 26.340 35.790 ;
        RECT 27.340 34.790 28.340 35.790 ;
        RECT 29.340 34.790 30.340 35.790 ;
        RECT 31.340 34.790 32.340 35.790 ;
        RECT 33.340 34.790 34.340 35.790 ;
        RECT 35.340 34.790 36.340 35.790 ;
        RECT 37.340 34.790 38.340 35.790 ;
        RECT 39.340 34.790 40.340 35.790 ;
        RECT 41.340 34.790 42.340 35.790 ;
        RECT 43.340 34.790 44.340 35.790 ;
        RECT 45.340 34.790 46.340 35.790 ;
        RECT 47.340 34.790 48.340 35.790 ;
        RECT 49.340 34.790 50.340 35.790 ;
        RECT 51.340 34.790 52.340 35.790 ;
        RECT 53.340 34.790 54.340 35.790 ;
        RECT 55.340 34.790 56.340 35.790 ;
        RECT 57.340 34.790 58.340 35.790 ;
        RECT 59.340 34.790 60.340 35.790 ;
        RECT 61.340 34.790 62.340 35.790 ;
        RECT 63.340 34.790 64.340 35.790 ;
        RECT 65.340 34.790 66.340 35.790 ;
        RECT 67.340 34.790 68.340 35.790 ;
        RECT 69.340 34.790 70.340 35.790 ;
        RECT 71.340 34.790 72.340 35.790 ;
        RECT 73.340 34.790 74.340 35.790 ;
        RECT 86.775 34.790 87.775 35.790 ;
        RECT 88.775 34.790 89.775 35.790 ;
        RECT 90.775 34.790 91.775 35.790 ;
        RECT 92.775 34.790 93.775 35.790 ;
        RECT 94.775 34.790 95.775 35.790 ;
        RECT 96.775 34.790 97.775 35.790 ;
        RECT 98.775 34.790 99.775 35.790 ;
        RECT 100.775 34.790 101.775 35.790 ;
        RECT 102.775 34.790 103.775 35.790 ;
        RECT 104.775 34.790 105.775 35.790 ;
        RECT 106.775 34.790 107.775 35.790 ;
        RECT 108.775 34.790 109.775 35.790 ;
        RECT 110.775 34.790 111.775 35.790 ;
        RECT 112.775 34.790 113.775 35.790 ;
        RECT 114.775 34.790 115.775 35.790 ;
        RECT 116.775 34.790 117.775 35.790 ;
        RECT 118.775 34.790 119.775 35.790 ;
        RECT 120.775 34.790 121.775 35.790 ;
        RECT 122.775 34.790 123.775 35.790 ;
        RECT 124.775 34.790 125.775 35.790 ;
        RECT 126.775 34.790 127.775 35.790 ;
        RECT 128.775 34.790 129.775 35.790 ;
        RECT 130.775 34.790 131.775 35.790 ;
        RECT 132.775 34.790 133.775 35.790 ;
        RECT 134.775 34.790 135.775 35.790 ;
        RECT 136.775 34.790 137.775 35.790 ;
        RECT 138.775 34.790 139.775 35.790 ;
        RECT 140.775 34.790 141.775 35.790 ;
        RECT 142.775 34.790 143.775 35.790 ;
        RECT 144.775 34.790 145.775 35.790 ;
        RECT 146.775 34.790 147.775 35.790 ;
        RECT 148.775 34.790 149.775 35.790 ;
        RECT 150.775 34.790 151.775 35.790 ;
        RECT 152.775 34.790 153.775 35.790 ;
        RECT 7.690 33.940 7.990 34.790 ;
        RECT 9.690 33.940 9.990 34.790 ;
        RECT 11.690 33.940 11.990 34.790 ;
        RECT 13.690 33.940 13.990 34.790 ;
        RECT 15.690 33.940 15.990 34.790 ;
        RECT 17.690 33.940 17.990 34.790 ;
        RECT 19.690 33.940 19.990 34.790 ;
        RECT 21.690 33.940 21.990 34.790 ;
        RECT 23.690 33.940 23.990 34.790 ;
        RECT 25.690 33.940 25.990 34.790 ;
        RECT 27.690 33.940 27.990 34.790 ;
        RECT 29.690 33.940 29.990 34.790 ;
        RECT 31.690 33.940 31.990 34.790 ;
        RECT 33.690 33.940 33.990 34.790 ;
        RECT 35.690 33.940 35.990 34.790 ;
        RECT 37.690 33.940 37.990 34.790 ;
        RECT 39.690 33.940 39.990 34.790 ;
        RECT 41.690 33.940 41.990 34.790 ;
        RECT 43.690 33.940 43.990 34.790 ;
        RECT 45.690 33.940 45.990 34.790 ;
        RECT 47.690 33.940 47.990 34.790 ;
        RECT 49.690 33.940 49.990 34.790 ;
        RECT 51.690 33.940 51.990 34.790 ;
        RECT 53.690 33.940 53.990 34.790 ;
        RECT 55.690 33.940 55.990 34.790 ;
        RECT 57.690 33.940 57.990 34.790 ;
        RECT 59.690 33.940 59.990 34.790 ;
        RECT 61.690 33.940 61.990 34.790 ;
        RECT 63.690 33.940 63.990 34.790 ;
        RECT 65.690 33.940 65.990 34.790 ;
        RECT 67.690 33.940 67.990 34.790 ;
        RECT 69.690 33.940 69.990 34.790 ;
        RECT 71.690 33.940 71.990 34.790 ;
        RECT 73.690 33.940 73.990 34.790 ;
        RECT 87.125 33.940 87.425 34.790 ;
        RECT 89.125 33.940 89.425 34.790 ;
        RECT 91.125 33.940 91.425 34.790 ;
        RECT 93.125 33.940 93.425 34.790 ;
        RECT 95.125 33.940 95.425 34.790 ;
        RECT 97.125 33.940 97.425 34.790 ;
        RECT 99.125 33.940 99.425 34.790 ;
        RECT 101.125 33.940 101.425 34.790 ;
        RECT 103.125 33.940 103.425 34.790 ;
        RECT 105.125 33.940 105.425 34.790 ;
        RECT 107.125 33.940 107.425 34.790 ;
        RECT 109.125 33.940 109.425 34.790 ;
        RECT 111.125 33.940 111.425 34.790 ;
        RECT 113.125 33.940 113.425 34.790 ;
        RECT 115.125 33.940 115.425 34.790 ;
        RECT 117.125 33.940 117.425 34.790 ;
        RECT 119.125 33.940 119.425 34.790 ;
        RECT 121.125 33.940 121.425 34.790 ;
        RECT 123.125 33.940 123.425 34.790 ;
        RECT 125.125 33.940 125.425 34.790 ;
        RECT 127.125 33.940 127.425 34.790 ;
        RECT 129.125 33.940 129.425 34.790 ;
        RECT 131.125 33.940 131.425 34.790 ;
        RECT 133.125 33.940 133.425 34.790 ;
        RECT 135.125 33.940 135.425 34.790 ;
        RECT 137.125 33.940 137.425 34.790 ;
        RECT 139.125 33.940 139.425 34.790 ;
        RECT 141.125 33.940 141.425 34.790 ;
        RECT 143.125 33.940 143.425 34.790 ;
        RECT 145.125 33.940 145.425 34.790 ;
        RECT 147.125 33.940 147.425 34.790 ;
        RECT 149.125 33.940 149.425 34.790 ;
        RECT 151.125 33.940 151.425 34.790 ;
        RECT 153.125 33.940 153.425 34.790 ;
        RECT 7.340 32.940 8.340 33.940 ;
        RECT 9.340 32.940 10.340 33.940 ;
        RECT 11.340 32.940 12.340 33.940 ;
        RECT 13.340 32.940 14.340 33.940 ;
        RECT 15.340 32.940 16.340 33.940 ;
        RECT 17.340 32.940 18.340 33.940 ;
        RECT 19.340 32.940 20.340 33.940 ;
        RECT 21.340 32.940 22.340 33.940 ;
        RECT 23.340 32.940 24.340 33.940 ;
        RECT 25.340 32.940 26.340 33.940 ;
        RECT 27.340 32.940 28.340 33.940 ;
        RECT 29.340 32.940 30.340 33.940 ;
        RECT 31.340 32.940 32.340 33.940 ;
        RECT 33.340 32.940 34.340 33.940 ;
        RECT 35.340 32.940 36.340 33.940 ;
        RECT 37.340 32.940 38.340 33.940 ;
        RECT 39.340 32.940 40.340 33.940 ;
        RECT 41.340 32.940 42.340 33.940 ;
        RECT 43.340 32.940 44.340 33.940 ;
        RECT 45.340 32.940 46.340 33.940 ;
        RECT 47.340 32.940 48.340 33.940 ;
        RECT 49.340 32.940 50.340 33.940 ;
        RECT 51.340 32.940 52.340 33.940 ;
        RECT 53.340 32.940 54.340 33.940 ;
        RECT 55.340 32.940 56.340 33.940 ;
        RECT 57.340 32.940 58.340 33.940 ;
        RECT 59.340 32.940 60.340 33.940 ;
        RECT 61.340 32.940 62.340 33.940 ;
        RECT 63.340 32.940 64.340 33.940 ;
        RECT 65.340 32.940 66.340 33.940 ;
        RECT 67.340 32.940 68.340 33.940 ;
        RECT 69.340 32.940 70.340 33.940 ;
        RECT 71.340 32.940 72.340 33.940 ;
        RECT 73.340 32.940 74.340 33.940 ;
        RECT 86.775 32.940 87.775 33.940 ;
        RECT 88.775 32.940 89.775 33.940 ;
        RECT 90.775 32.940 91.775 33.940 ;
        RECT 92.775 32.940 93.775 33.940 ;
        RECT 94.775 32.940 95.775 33.940 ;
        RECT 96.775 32.940 97.775 33.940 ;
        RECT 98.775 32.940 99.775 33.940 ;
        RECT 100.775 32.940 101.775 33.940 ;
        RECT 102.775 32.940 103.775 33.940 ;
        RECT 104.775 32.940 105.775 33.940 ;
        RECT 106.775 32.940 107.775 33.940 ;
        RECT 108.775 32.940 109.775 33.940 ;
        RECT 110.775 32.940 111.775 33.940 ;
        RECT 112.775 32.940 113.775 33.940 ;
        RECT 114.775 32.940 115.775 33.940 ;
        RECT 116.775 32.940 117.775 33.940 ;
        RECT 118.775 32.940 119.775 33.940 ;
        RECT 120.775 32.940 121.775 33.940 ;
        RECT 122.775 32.940 123.775 33.940 ;
        RECT 124.775 32.940 125.775 33.940 ;
        RECT 126.775 32.940 127.775 33.940 ;
        RECT 128.775 32.940 129.775 33.940 ;
        RECT 130.775 32.940 131.775 33.940 ;
        RECT 132.775 32.940 133.775 33.940 ;
        RECT 134.775 32.940 135.775 33.940 ;
        RECT 136.775 32.940 137.775 33.940 ;
        RECT 138.775 32.940 139.775 33.940 ;
        RECT 140.775 32.940 141.775 33.940 ;
        RECT 142.775 32.940 143.775 33.940 ;
        RECT 144.775 32.940 145.775 33.940 ;
        RECT 146.775 32.940 147.775 33.940 ;
        RECT 148.775 32.940 149.775 33.940 ;
        RECT 150.775 32.940 151.775 33.940 ;
        RECT 152.775 32.940 153.775 33.940 ;
        RECT 7.690 32.090 7.990 32.940 ;
        RECT 9.690 32.090 9.990 32.940 ;
        RECT 11.690 32.090 11.990 32.940 ;
        RECT 13.690 32.090 13.990 32.940 ;
        RECT 15.690 32.090 15.990 32.940 ;
        RECT 17.690 32.090 17.990 32.940 ;
        RECT 19.690 32.090 19.990 32.940 ;
        RECT 21.690 32.090 21.990 32.940 ;
        RECT 23.690 32.090 23.990 32.940 ;
        RECT 25.690 32.090 25.990 32.940 ;
        RECT 27.690 32.090 27.990 32.940 ;
        RECT 29.690 32.090 29.990 32.940 ;
        RECT 31.690 32.090 31.990 32.940 ;
        RECT 33.690 32.090 33.990 32.940 ;
        RECT 35.690 32.090 35.990 32.940 ;
        RECT 37.690 32.090 37.990 32.940 ;
        RECT 39.690 32.090 39.990 32.940 ;
        RECT 41.690 32.090 41.990 32.940 ;
        RECT 43.690 32.090 43.990 32.940 ;
        RECT 45.690 32.090 45.990 32.940 ;
        RECT 47.690 32.090 47.990 32.940 ;
        RECT 49.690 32.090 49.990 32.940 ;
        RECT 51.690 32.090 51.990 32.940 ;
        RECT 53.690 32.090 53.990 32.940 ;
        RECT 55.690 32.090 55.990 32.940 ;
        RECT 57.690 32.090 57.990 32.940 ;
        RECT 59.690 32.090 59.990 32.940 ;
        RECT 61.690 32.090 61.990 32.940 ;
        RECT 63.690 32.090 63.990 32.940 ;
        RECT 65.690 32.090 65.990 32.940 ;
        RECT 67.690 32.090 67.990 32.940 ;
        RECT 69.690 32.090 69.990 32.940 ;
        RECT 71.690 32.090 71.990 32.940 ;
        RECT 73.690 32.090 73.990 32.940 ;
        RECT 87.125 32.090 87.425 32.940 ;
        RECT 89.125 32.090 89.425 32.940 ;
        RECT 91.125 32.090 91.425 32.940 ;
        RECT 93.125 32.090 93.425 32.940 ;
        RECT 95.125 32.090 95.425 32.940 ;
        RECT 97.125 32.090 97.425 32.940 ;
        RECT 99.125 32.090 99.425 32.940 ;
        RECT 101.125 32.090 101.425 32.940 ;
        RECT 103.125 32.090 103.425 32.940 ;
        RECT 105.125 32.090 105.425 32.940 ;
        RECT 107.125 32.090 107.425 32.940 ;
        RECT 109.125 32.090 109.425 32.940 ;
        RECT 111.125 32.090 111.425 32.940 ;
        RECT 113.125 32.090 113.425 32.940 ;
        RECT 115.125 32.090 115.425 32.940 ;
        RECT 117.125 32.090 117.425 32.940 ;
        RECT 119.125 32.090 119.425 32.940 ;
        RECT 121.125 32.090 121.425 32.940 ;
        RECT 123.125 32.090 123.425 32.940 ;
        RECT 125.125 32.090 125.425 32.940 ;
        RECT 127.125 32.090 127.425 32.940 ;
        RECT 129.125 32.090 129.425 32.940 ;
        RECT 131.125 32.090 131.425 32.940 ;
        RECT 133.125 32.090 133.425 32.940 ;
        RECT 135.125 32.090 135.425 32.940 ;
        RECT 137.125 32.090 137.425 32.940 ;
        RECT 139.125 32.090 139.425 32.940 ;
        RECT 141.125 32.090 141.425 32.940 ;
        RECT 143.125 32.090 143.425 32.940 ;
        RECT 145.125 32.090 145.425 32.940 ;
        RECT 147.125 32.090 147.425 32.940 ;
        RECT 149.125 32.090 149.425 32.940 ;
        RECT 151.125 32.090 151.425 32.940 ;
        RECT 153.125 32.090 153.425 32.940 ;
        RECT 7.340 31.090 8.340 32.090 ;
        RECT 9.340 31.090 10.340 32.090 ;
        RECT 11.340 31.090 12.340 32.090 ;
        RECT 13.340 31.090 14.340 32.090 ;
        RECT 15.340 31.090 16.340 32.090 ;
        RECT 17.340 31.090 18.340 32.090 ;
        RECT 19.340 31.090 20.340 32.090 ;
        RECT 21.340 31.090 22.340 32.090 ;
        RECT 23.340 31.090 24.340 32.090 ;
        RECT 25.340 31.090 26.340 32.090 ;
        RECT 27.340 31.090 28.340 32.090 ;
        RECT 29.340 31.090 30.340 32.090 ;
        RECT 31.340 31.090 32.340 32.090 ;
        RECT 33.340 31.090 34.340 32.090 ;
        RECT 35.340 31.090 36.340 32.090 ;
        RECT 37.340 31.090 38.340 32.090 ;
        RECT 39.340 31.090 40.340 32.090 ;
        RECT 41.340 31.090 42.340 32.090 ;
        RECT 43.340 31.090 44.340 32.090 ;
        RECT 45.340 31.090 46.340 32.090 ;
        RECT 47.340 31.090 48.340 32.090 ;
        RECT 49.340 31.090 50.340 32.090 ;
        RECT 51.340 31.090 52.340 32.090 ;
        RECT 53.340 31.090 54.340 32.090 ;
        RECT 55.340 31.090 56.340 32.090 ;
        RECT 57.340 31.090 58.340 32.090 ;
        RECT 59.340 31.090 60.340 32.090 ;
        RECT 61.340 31.090 62.340 32.090 ;
        RECT 63.340 31.090 64.340 32.090 ;
        RECT 65.340 31.090 66.340 32.090 ;
        RECT 67.340 31.090 68.340 32.090 ;
        RECT 69.340 31.090 70.340 32.090 ;
        RECT 71.340 31.090 72.340 32.090 ;
        RECT 73.340 31.090 74.340 32.090 ;
        RECT 86.775 31.090 87.775 32.090 ;
        RECT 88.775 31.090 89.775 32.090 ;
        RECT 90.775 31.090 91.775 32.090 ;
        RECT 92.775 31.090 93.775 32.090 ;
        RECT 94.775 31.090 95.775 32.090 ;
        RECT 96.775 31.090 97.775 32.090 ;
        RECT 98.775 31.090 99.775 32.090 ;
        RECT 100.775 31.090 101.775 32.090 ;
        RECT 102.775 31.090 103.775 32.090 ;
        RECT 104.775 31.090 105.775 32.090 ;
        RECT 106.775 31.090 107.775 32.090 ;
        RECT 108.775 31.090 109.775 32.090 ;
        RECT 110.775 31.090 111.775 32.090 ;
        RECT 112.775 31.090 113.775 32.090 ;
        RECT 114.775 31.090 115.775 32.090 ;
        RECT 116.775 31.090 117.775 32.090 ;
        RECT 118.775 31.090 119.775 32.090 ;
        RECT 120.775 31.090 121.775 32.090 ;
        RECT 122.775 31.090 123.775 32.090 ;
        RECT 124.775 31.090 125.775 32.090 ;
        RECT 126.775 31.090 127.775 32.090 ;
        RECT 128.775 31.090 129.775 32.090 ;
        RECT 130.775 31.090 131.775 32.090 ;
        RECT 132.775 31.090 133.775 32.090 ;
        RECT 134.775 31.090 135.775 32.090 ;
        RECT 136.775 31.090 137.775 32.090 ;
        RECT 138.775 31.090 139.775 32.090 ;
        RECT 140.775 31.090 141.775 32.090 ;
        RECT 142.775 31.090 143.775 32.090 ;
        RECT 144.775 31.090 145.775 32.090 ;
        RECT 146.775 31.090 147.775 32.090 ;
        RECT 148.775 31.090 149.775 32.090 ;
        RECT 150.775 31.090 151.775 32.090 ;
        RECT 152.775 31.090 153.775 32.090 ;
        RECT 7.690 30.240 7.990 31.090 ;
        RECT 9.690 30.240 9.990 31.090 ;
        RECT 11.690 30.240 11.990 31.090 ;
        RECT 13.690 30.240 13.990 31.090 ;
        RECT 15.690 30.240 15.990 31.090 ;
        RECT 17.690 30.240 17.990 31.090 ;
        RECT 19.690 30.240 19.990 31.090 ;
        RECT 21.690 30.240 21.990 31.090 ;
        RECT 23.690 30.240 23.990 31.090 ;
        RECT 25.690 30.240 25.990 31.090 ;
        RECT 27.690 30.240 27.990 31.090 ;
        RECT 29.690 30.240 29.990 31.090 ;
        RECT 31.690 30.240 31.990 31.090 ;
        RECT 33.690 30.240 33.990 31.090 ;
        RECT 35.690 30.240 35.990 31.090 ;
        RECT 37.690 30.240 37.990 31.090 ;
        RECT 39.690 30.240 39.990 31.090 ;
        RECT 41.690 30.240 41.990 31.090 ;
        RECT 43.690 30.240 43.990 31.090 ;
        RECT 45.690 30.240 45.990 31.090 ;
        RECT 47.690 30.240 47.990 31.090 ;
        RECT 49.690 30.240 49.990 31.090 ;
        RECT 51.690 30.240 51.990 31.090 ;
        RECT 53.690 30.240 53.990 31.090 ;
        RECT 55.690 30.240 55.990 31.090 ;
        RECT 57.690 30.240 57.990 31.090 ;
        RECT 59.690 30.240 59.990 31.090 ;
        RECT 61.690 30.240 61.990 31.090 ;
        RECT 63.690 30.240 63.990 31.090 ;
        RECT 65.690 30.240 65.990 31.090 ;
        RECT 67.690 30.240 67.990 31.090 ;
        RECT 69.690 30.240 69.990 31.090 ;
        RECT 71.690 30.240 71.990 31.090 ;
        RECT 73.690 30.240 73.990 31.090 ;
        RECT 87.125 30.240 87.425 31.090 ;
        RECT 89.125 30.240 89.425 31.090 ;
        RECT 91.125 30.240 91.425 31.090 ;
        RECT 93.125 30.240 93.425 31.090 ;
        RECT 95.125 30.240 95.425 31.090 ;
        RECT 97.125 30.240 97.425 31.090 ;
        RECT 99.125 30.240 99.425 31.090 ;
        RECT 101.125 30.240 101.425 31.090 ;
        RECT 103.125 30.240 103.425 31.090 ;
        RECT 105.125 30.240 105.425 31.090 ;
        RECT 107.125 30.240 107.425 31.090 ;
        RECT 109.125 30.240 109.425 31.090 ;
        RECT 111.125 30.240 111.425 31.090 ;
        RECT 113.125 30.240 113.425 31.090 ;
        RECT 115.125 30.240 115.425 31.090 ;
        RECT 117.125 30.240 117.425 31.090 ;
        RECT 119.125 30.240 119.425 31.090 ;
        RECT 121.125 30.240 121.425 31.090 ;
        RECT 123.125 30.240 123.425 31.090 ;
        RECT 125.125 30.240 125.425 31.090 ;
        RECT 127.125 30.240 127.425 31.090 ;
        RECT 129.125 30.240 129.425 31.090 ;
        RECT 131.125 30.240 131.425 31.090 ;
        RECT 133.125 30.240 133.425 31.090 ;
        RECT 135.125 30.240 135.425 31.090 ;
        RECT 137.125 30.240 137.425 31.090 ;
        RECT 139.125 30.240 139.425 31.090 ;
        RECT 141.125 30.240 141.425 31.090 ;
        RECT 143.125 30.240 143.425 31.090 ;
        RECT 145.125 30.240 145.425 31.090 ;
        RECT 147.125 30.240 147.425 31.090 ;
        RECT 149.125 30.240 149.425 31.090 ;
        RECT 151.125 30.240 151.425 31.090 ;
        RECT 153.125 30.240 153.425 31.090 ;
        RECT 7.340 29.240 8.340 30.240 ;
        RECT 9.340 29.240 10.340 30.240 ;
        RECT 11.340 29.240 12.340 30.240 ;
        RECT 13.340 29.240 14.340 30.240 ;
        RECT 15.340 29.240 16.340 30.240 ;
        RECT 17.340 29.240 18.340 30.240 ;
        RECT 19.340 29.240 20.340 30.240 ;
        RECT 21.340 29.240 22.340 30.240 ;
        RECT 23.340 29.240 24.340 30.240 ;
        RECT 25.340 29.240 26.340 30.240 ;
        RECT 27.340 29.240 28.340 30.240 ;
        RECT 29.340 29.240 30.340 30.240 ;
        RECT 31.340 29.240 32.340 30.240 ;
        RECT 33.340 29.240 34.340 30.240 ;
        RECT 35.340 29.240 36.340 30.240 ;
        RECT 37.340 29.240 38.340 30.240 ;
        RECT 39.340 29.240 40.340 30.240 ;
        RECT 41.340 29.240 42.340 30.240 ;
        RECT 43.340 29.240 44.340 30.240 ;
        RECT 45.340 29.240 46.340 30.240 ;
        RECT 47.340 29.240 48.340 30.240 ;
        RECT 49.340 29.240 50.340 30.240 ;
        RECT 51.340 29.240 52.340 30.240 ;
        RECT 53.340 29.240 54.340 30.240 ;
        RECT 55.340 29.240 56.340 30.240 ;
        RECT 57.340 29.240 58.340 30.240 ;
        RECT 59.340 29.240 60.340 30.240 ;
        RECT 61.340 29.240 62.340 30.240 ;
        RECT 63.340 29.240 64.340 30.240 ;
        RECT 65.340 29.240 66.340 30.240 ;
        RECT 67.340 29.240 68.340 30.240 ;
        RECT 69.340 29.240 70.340 30.240 ;
        RECT 71.340 29.240 72.340 30.240 ;
        RECT 73.340 29.240 74.340 30.240 ;
        RECT 86.775 29.240 87.775 30.240 ;
        RECT 88.775 29.240 89.775 30.240 ;
        RECT 90.775 29.240 91.775 30.240 ;
        RECT 92.775 29.240 93.775 30.240 ;
        RECT 94.775 29.240 95.775 30.240 ;
        RECT 96.775 29.240 97.775 30.240 ;
        RECT 98.775 29.240 99.775 30.240 ;
        RECT 100.775 29.240 101.775 30.240 ;
        RECT 102.775 29.240 103.775 30.240 ;
        RECT 104.775 29.240 105.775 30.240 ;
        RECT 106.775 29.240 107.775 30.240 ;
        RECT 108.775 29.240 109.775 30.240 ;
        RECT 110.775 29.240 111.775 30.240 ;
        RECT 112.775 29.240 113.775 30.240 ;
        RECT 114.775 29.240 115.775 30.240 ;
        RECT 116.775 29.240 117.775 30.240 ;
        RECT 118.775 29.240 119.775 30.240 ;
        RECT 120.775 29.240 121.775 30.240 ;
        RECT 122.775 29.240 123.775 30.240 ;
        RECT 124.775 29.240 125.775 30.240 ;
        RECT 126.775 29.240 127.775 30.240 ;
        RECT 128.775 29.240 129.775 30.240 ;
        RECT 130.775 29.240 131.775 30.240 ;
        RECT 132.775 29.240 133.775 30.240 ;
        RECT 134.775 29.240 135.775 30.240 ;
        RECT 136.775 29.240 137.775 30.240 ;
        RECT 138.775 29.240 139.775 30.240 ;
        RECT 140.775 29.240 141.775 30.240 ;
        RECT 142.775 29.240 143.775 30.240 ;
        RECT 144.775 29.240 145.775 30.240 ;
        RECT 146.775 29.240 147.775 30.240 ;
        RECT 148.775 29.240 149.775 30.240 ;
        RECT 150.775 29.240 151.775 30.240 ;
        RECT 152.775 29.240 153.775 30.240 ;
        RECT 7.690 28.390 7.990 29.240 ;
        RECT 9.690 28.390 9.990 29.240 ;
        RECT 11.690 28.390 11.990 29.240 ;
        RECT 13.690 28.390 13.990 29.240 ;
        RECT 15.690 28.390 15.990 29.240 ;
        RECT 17.690 28.390 17.990 29.240 ;
        RECT 19.690 28.390 19.990 29.240 ;
        RECT 21.690 28.390 21.990 29.240 ;
        RECT 23.690 28.390 23.990 29.240 ;
        RECT 25.690 28.390 25.990 29.240 ;
        RECT 27.690 28.390 27.990 29.240 ;
        RECT 29.690 28.390 29.990 29.240 ;
        RECT 31.690 28.390 31.990 29.240 ;
        RECT 33.690 28.390 33.990 29.240 ;
        RECT 35.690 28.390 35.990 29.240 ;
        RECT 37.690 28.390 37.990 29.240 ;
        RECT 39.690 28.390 39.990 29.240 ;
        RECT 41.690 28.390 41.990 29.240 ;
        RECT 43.690 28.390 43.990 29.240 ;
        RECT 45.690 28.390 45.990 29.240 ;
        RECT 47.690 28.390 47.990 29.240 ;
        RECT 49.690 28.390 49.990 29.240 ;
        RECT 51.690 28.390 51.990 29.240 ;
        RECT 53.690 28.390 53.990 29.240 ;
        RECT 55.690 28.390 55.990 29.240 ;
        RECT 57.690 28.390 57.990 29.240 ;
        RECT 59.690 28.390 59.990 29.240 ;
        RECT 61.690 28.390 61.990 29.240 ;
        RECT 63.690 28.390 63.990 29.240 ;
        RECT 65.690 28.390 65.990 29.240 ;
        RECT 67.690 28.390 67.990 29.240 ;
        RECT 69.690 28.390 69.990 29.240 ;
        RECT 71.690 28.390 71.990 29.240 ;
        RECT 73.690 28.390 73.990 29.240 ;
        RECT 87.125 28.390 87.425 29.240 ;
        RECT 89.125 28.390 89.425 29.240 ;
        RECT 91.125 28.390 91.425 29.240 ;
        RECT 93.125 28.390 93.425 29.240 ;
        RECT 95.125 28.390 95.425 29.240 ;
        RECT 97.125 28.390 97.425 29.240 ;
        RECT 99.125 28.390 99.425 29.240 ;
        RECT 101.125 28.390 101.425 29.240 ;
        RECT 103.125 28.390 103.425 29.240 ;
        RECT 105.125 28.390 105.425 29.240 ;
        RECT 107.125 28.390 107.425 29.240 ;
        RECT 109.125 28.390 109.425 29.240 ;
        RECT 111.125 28.390 111.425 29.240 ;
        RECT 113.125 28.390 113.425 29.240 ;
        RECT 115.125 28.390 115.425 29.240 ;
        RECT 117.125 28.390 117.425 29.240 ;
        RECT 119.125 28.390 119.425 29.240 ;
        RECT 121.125 28.390 121.425 29.240 ;
        RECT 123.125 28.390 123.425 29.240 ;
        RECT 125.125 28.390 125.425 29.240 ;
        RECT 127.125 28.390 127.425 29.240 ;
        RECT 129.125 28.390 129.425 29.240 ;
        RECT 131.125 28.390 131.425 29.240 ;
        RECT 133.125 28.390 133.425 29.240 ;
        RECT 135.125 28.390 135.425 29.240 ;
        RECT 137.125 28.390 137.425 29.240 ;
        RECT 139.125 28.390 139.425 29.240 ;
        RECT 141.125 28.390 141.425 29.240 ;
        RECT 143.125 28.390 143.425 29.240 ;
        RECT 145.125 28.390 145.425 29.240 ;
        RECT 147.125 28.390 147.425 29.240 ;
        RECT 149.125 28.390 149.425 29.240 ;
        RECT 151.125 28.390 151.425 29.240 ;
        RECT 153.125 28.390 153.425 29.240 ;
        RECT 7.340 27.390 8.340 28.390 ;
        RECT 9.340 27.390 10.340 28.390 ;
        RECT 11.340 27.390 12.340 28.390 ;
        RECT 13.340 27.390 14.340 28.390 ;
        RECT 15.340 27.390 16.340 28.390 ;
        RECT 17.340 27.390 18.340 28.390 ;
        RECT 19.340 27.390 20.340 28.390 ;
        RECT 21.340 27.390 22.340 28.390 ;
        RECT 23.340 27.390 24.340 28.390 ;
        RECT 25.340 27.390 26.340 28.390 ;
        RECT 27.340 27.390 28.340 28.390 ;
        RECT 29.340 27.390 30.340 28.390 ;
        RECT 31.340 27.390 32.340 28.390 ;
        RECT 33.340 27.390 34.340 28.390 ;
        RECT 35.340 27.390 36.340 28.390 ;
        RECT 37.340 27.390 38.340 28.390 ;
        RECT 39.340 27.390 40.340 28.390 ;
        RECT 41.340 27.390 42.340 28.390 ;
        RECT 43.340 27.390 44.340 28.390 ;
        RECT 45.340 27.390 46.340 28.390 ;
        RECT 47.340 27.390 48.340 28.390 ;
        RECT 49.340 27.390 50.340 28.390 ;
        RECT 51.340 27.390 52.340 28.390 ;
        RECT 53.340 27.390 54.340 28.390 ;
        RECT 55.340 27.390 56.340 28.390 ;
        RECT 57.340 27.390 58.340 28.390 ;
        RECT 59.340 27.390 60.340 28.390 ;
        RECT 61.340 27.390 62.340 28.390 ;
        RECT 63.340 27.390 64.340 28.390 ;
        RECT 65.340 27.390 66.340 28.390 ;
        RECT 67.340 27.390 68.340 28.390 ;
        RECT 69.340 27.390 70.340 28.390 ;
        RECT 71.340 27.390 72.340 28.390 ;
        RECT 73.340 27.390 74.340 28.390 ;
        RECT 86.775 27.390 87.775 28.390 ;
        RECT 88.775 27.390 89.775 28.390 ;
        RECT 90.775 27.390 91.775 28.390 ;
        RECT 92.775 27.390 93.775 28.390 ;
        RECT 94.775 27.390 95.775 28.390 ;
        RECT 96.775 27.390 97.775 28.390 ;
        RECT 98.775 27.390 99.775 28.390 ;
        RECT 100.775 27.390 101.775 28.390 ;
        RECT 102.775 27.390 103.775 28.390 ;
        RECT 104.775 27.390 105.775 28.390 ;
        RECT 106.775 27.390 107.775 28.390 ;
        RECT 108.775 27.390 109.775 28.390 ;
        RECT 110.775 27.390 111.775 28.390 ;
        RECT 112.775 27.390 113.775 28.390 ;
        RECT 114.775 27.390 115.775 28.390 ;
        RECT 116.775 27.390 117.775 28.390 ;
        RECT 118.775 27.390 119.775 28.390 ;
        RECT 120.775 27.390 121.775 28.390 ;
        RECT 122.775 27.390 123.775 28.390 ;
        RECT 124.775 27.390 125.775 28.390 ;
        RECT 126.775 27.390 127.775 28.390 ;
        RECT 128.775 27.390 129.775 28.390 ;
        RECT 130.775 27.390 131.775 28.390 ;
        RECT 132.775 27.390 133.775 28.390 ;
        RECT 134.775 27.390 135.775 28.390 ;
        RECT 136.775 27.390 137.775 28.390 ;
        RECT 138.775 27.390 139.775 28.390 ;
        RECT 140.775 27.390 141.775 28.390 ;
        RECT 142.775 27.390 143.775 28.390 ;
        RECT 144.775 27.390 145.775 28.390 ;
        RECT 146.775 27.390 147.775 28.390 ;
        RECT 148.775 27.390 149.775 28.390 ;
        RECT 150.775 27.390 151.775 28.390 ;
        RECT 152.775 27.390 153.775 28.390 ;
        RECT 7.690 26.540 7.990 27.390 ;
        RECT 9.690 26.540 9.990 27.390 ;
        RECT 11.690 26.540 11.990 27.390 ;
        RECT 13.690 26.540 13.990 27.390 ;
        RECT 15.690 26.540 15.990 27.390 ;
        RECT 17.690 26.540 17.990 27.390 ;
        RECT 19.690 26.540 19.990 27.390 ;
        RECT 21.690 26.540 21.990 27.390 ;
        RECT 23.690 26.540 23.990 27.390 ;
        RECT 25.690 26.540 25.990 27.390 ;
        RECT 27.690 26.540 27.990 27.390 ;
        RECT 29.690 26.540 29.990 27.390 ;
        RECT 31.690 26.540 31.990 27.390 ;
        RECT 33.690 26.540 33.990 27.390 ;
        RECT 35.690 26.540 35.990 27.390 ;
        RECT 37.690 26.540 37.990 27.390 ;
        RECT 39.690 26.540 39.990 27.390 ;
        RECT 41.690 26.540 41.990 27.390 ;
        RECT 43.690 26.540 43.990 27.390 ;
        RECT 45.690 26.540 45.990 27.390 ;
        RECT 47.690 26.540 47.990 27.390 ;
        RECT 49.690 26.540 49.990 27.390 ;
        RECT 51.690 26.540 51.990 27.390 ;
        RECT 53.690 26.540 53.990 27.390 ;
        RECT 55.690 26.540 55.990 27.390 ;
        RECT 57.690 26.540 57.990 27.390 ;
        RECT 59.690 26.540 59.990 27.390 ;
        RECT 61.690 26.540 61.990 27.390 ;
        RECT 63.690 26.540 63.990 27.390 ;
        RECT 65.690 26.540 65.990 27.390 ;
        RECT 67.690 26.540 67.990 27.390 ;
        RECT 69.690 26.540 69.990 27.390 ;
        RECT 71.690 26.540 71.990 27.390 ;
        RECT 73.690 26.540 73.990 27.390 ;
        RECT 87.125 26.540 87.425 27.390 ;
        RECT 89.125 26.540 89.425 27.390 ;
        RECT 91.125 26.540 91.425 27.390 ;
        RECT 93.125 26.540 93.425 27.390 ;
        RECT 95.125 26.540 95.425 27.390 ;
        RECT 97.125 26.540 97.425 27.390 ;
        RECT 99.125 26.540 99.425 27.390 ;
        RECT 101.125 26.540 101.425 27.390 ;
        RECT 103.125 26.540 103.425 27.390 ;
        RECT 105.125 26.540 105.425 27.390 ;
        RECT 107.125 26.540 107.425 27.390 ;
        RECT 109.125 26.540 109.425 27.390 ;
        RECT 111.125 26.540 111.425 27.390 ;
        RECT 113.125 26.540 113.425 27.390 ;
        RECT 115.125 26.540 115.425 27.390 ;
        RECT 117.125 26.540 117.425 27.390 ;
        RECT 119.125 26.540 119.425 27.390 ;
        RECT 121.125 26.540 121.425 27.390 ;
        RECT 123.125 26.540 123.425 27.390 ;
        RECT 125.125 26.540 125.425 27.390 ;
        RECT 127.125 26.540 127.425 27.390 ;
        RECT 129.125 26.540 129.425 27.390 ;
        RECT 131.125 26.540 131.425 27.390 ;
        RECT 133.125 26.540 133.425 27.390 ;
        RECT 135.125 26.540 135.425 27.390 ;
        RECT 137.125 26.540 137.425 27.390 ;
        RECT 139.125 26.540 139.425 27.390 ;
        RECT 141.125 26.540 141.425 27.390 ;
        RECT 143.125 26.540 143.425 27.390 ;
        RECT 145.125 26.540 145.425 27.390 ;
        RECT 147.125 26.540 147.425 27.390 ;
        RECT 149.125 26.540 149.425 27.390 ;
        RECT 151.125 26.540 151.425 27.390 ;
        RECT 153.125 26.540 153.425 27.390 ;
        RECT 7.340 25.540 8.340 26.540 ;
        RECT 9.340 25.540 10.340 26.540 ;
        RECT 11.340 25.540 12.340 26.540 ;
        RECT 13.340 25.540 14.340 26.540 ;
        RECT 15.340 25.540 16.340 26.540 ;
        RECT 17.340 25.540 18.340 26.540 ;
        RECT 19.340 25.540 20.340 26.540 ;
        RECT 21.340 25.540 22.340 26.540 ;
        RECT 23.340 25.540 24.340 26.540 ;
        RECT 25.340 25.540 26.340 26.540 ;
        RECT 27.340 25.540 28.340 26.540 ;
        RECT 29.340 25.540 30.340 26.540 ;
        RECT 31.340 25.540 32.340 26.540 ;
        RECT 33.340 25.540 34.340 26.540 ;
        RECT 35.340 25.540 36.340 26.540 ;
        RECT 37.340 25.540 38.340 26.540 ;
        RECT 39.340 25.540 40.340 26.540 ;
        RECT 41.340 25.540 42.340 26.540 ;
        RECT 43.340 25.540 44.340 26.540 ;
        RECT 45.340 25.540 46.340 26.540 ;
        RECT 47.340 25.540 48.340 26.540 ;
        RECT 49.340 25.540 50.340 26.540 ;
        RECT 51.340 25.540 52.340 26.540 ;
        RECT 53.340 25.540 54.340 26.540 ;
        RECT 55.340 25.540 56.340 26.540 ;
        RECT 57.340 25.540 58.340 26.540 ;
        RECT 59.340 25.540 60.340 26.540 ;
        RECT 61.340 25.540 62.340 26.540 ;
        RECT 63.340 25.540 64.340 26.540 ;
        RECT 65.340 25.540 66.340 26.540 ;
        RECT 67.340 25.540 68.340 26.540 ;
        RECT 69.340 25.540 70.340 26.540 ;
        RECT 71.340 25.540 72.340 26.540 ;
        RECT 73.340 25.540 74.340 26.540 ;
        RECT 86.775 25.540 87.775 26.540 ;
        RECT 88.775 25.540 89.775 26.540 ;
        RECT 90.775 25.540 91.775 26.540 ;
        RECT 92.775 25.540 93.775 26.540 ;
        RECT 94.775 25.540 95.775 26.540 ;
        RECT 96.775 25.540 97.775 26.540 ;
        RECT 98.775 25.540 99.775 26.540 ;
        RECT 100.775 25.540 101.775 26.540 ;
        RECT 102.775 25.540 103.775 26.540 ;
        RECT 104.775 25.540 105.775 26.540 ;
        RECT 106.775 25.540 107.775 26.540 ;
        RECT 108.775 25.540 109.775 26.540 ;
        RECT 110.775 25.540 111.775 26.540 ;
        RECT 112.775 25.540 113.775 26.540 ;
        RECT 114.775 25.540 115.775 26.540 ;
        RECT 116.775 25.540 117.775 26.540 ;
        RECT 118.775 25.540 119.775 26.540 ;
        RECT 120.775 25.540 121.775 26.540 ;
        RECT 122.775 25.540 123.775 26.540 ;
        RECT 124.775 25.540 125.775 26.540 ;
        RECT 126.775 25.540 127.775 26.540 ;
        RECT 128.775 25.540 129.775 26.540 ;
        RECT 130.775 25.540 131.775 26.540 ;
        RECT 132.775 25.540 133.775 26.540 ;
        RECT 134.775 25.540 135.775 26.540 ;
        RECT 136.775 25.540 137.775 26.540 ;
        RECT 138.775 25.540 139.775 26.540 ;
        RECT 140.775 25.540 141.775 26.540 ;
        RECT 142.775 25.540 143.775 26.540 ;
        RECT 144.775 25.540 145.775 26.540 ;
        RECT 146.775 25.540 147.775 26.540 ;
        RECT 148.775 25.540 149.775 26.540 ;
        RECT 150.775 25.540 151.775 26.540 ;
        RECT 152.775 25.540 153.775 26.540 ;
        RECT 7.690 24.690 7.990 25.540 ;
        RECT 9.690 24.690 9.990 25.540 ;
        RECT 11.690 24.690 11.990 25.540 ;
        RECT 13.690 24.690 13.990 25.540 ;
        RECT 15.690 24.690 15.990 25.540 ;
        RECT 17.690 24.690 17.990 25.540 ;
        RECT 19.690 24.690 19.990 25.540 ;
        RECT 21.690 24.690 21.990 25.540 ;
        RECT 23.690 24.690 23.990 25.540 ;
        RECT 25.690 24.690 25.990 25.540 ;
        RECT 27.690 24.690 27.990 25.540 ;
        RECT 29.690 24.690 29.990 25.540 ;
        RECT 31.690 24.690 31.990 25.540 ;
        RECT 33.690 24.690 33.990 25.540 ;
        RECT 35.690 24.690 35.990 25.540 ;
        RECT 37.690 24.690 37.990 25.540 ;
        RECT 39.690 24.690 39.990 25.540 ;
        RECT 41.690 24.690 41.990 25.540 ;
        RECT 43.690 24.690 43.990 25.540 ;
        RECT 45.690 24.690 45.990 25.540 ;
        RECT 47.690 24.690 47.990 25.540 ;
        RECT 49.690 24.690 49.990 25.540 ;
        RECT 51.690 24.690 51.990 25.540 ;
        RECT 53.690 24.690 53.990 25.540 ;
        RECT 55.690 24.690 55.990 25.540 ;
        RECT 57.690 24.690 57.990 25.540 ;
        RECT 59.690 24.690 59.990 25.540 ;
        RECT 61.690 24.690 61.990 25.540 ;
        RECT 63.690 24.690 63.990 25.540 ;
        RECT 65.690 24.690 65.990 25.540 ;
        RECT 67.690 24.690 67.990 25.540 ;
        RECT 69.690 24.690 69.990 25.540 ;
        RECT 71.690 24.690 71.990 25.540 ;
        RECT 73.690 24.690 73.990 25.540 ;
        RECT 87.125 24.690 87.425 25.540 ;
        RECT 89.125 24.690 89.425 25.540 ;
        RECT 91.125 24.690 91.425 25.540 ;
        RECT 93.125 24.690 93.425 25.540 ;
        RECT 95.125 24.690 95.425 25.540 ;
        RECT 97.125 24.690 97.425 25.540 ;
        RECT 99.125 24.690 99.425 25.540 ;
        RECT 101.125 24.690 101.425 25.540 ;
        RECT 103.125 24.690 103.425 25.540 ;
        RECT 105.125 24.690 105.425 25.540 ;
        RECT 107.125 24.690 107.425 25.540 ;
        RECT 109.125 24.690 109.425 25.540 ;
        RECT 111.125 24.690 111.425 25.540 ;
        RECT 113.125 24.690 113.425 25.540 ;
        RECT 115.125 24.690 115.425 25.540 ;
        RECT 117.125 24.690 117.425 25.540 ;
        RECT 119.125 24.690 119.425 25.540 ;
        RECT 121.125 24.690 121.425 25.540 ;
        RECT 123.125 24.690 123.425 25.540 ;
        RECT 125.125 24.690 125.425 25.540 ;
        RECT 127.125 24.690 127.425 25.540 ;
        RECT 129.125 24.690 129.425 25.540 ;
        RECT 131.125 24.690 131.425 25.540 ;
        RECT 133.125 24.690 133.425 25.540 ;
        RECT 135.125 24.690 135.425 25.540 ;
        RECT 137.125 24.690 137.425 25.540 ;
        RECT 139.125 24.690 139.425 25.540 ;
        RECT 141.125 24.690 141.425 25.540 ;
        RECT 143.125 24.690 143.425 25.540 ;
        RECT 145.125 24.690 145.425 25.540 ;
        RECT 147.125 24.690 147.425 25.540 ;
        RECT 149.125 24.690 149.425 25.540 ;
        RECT 151.125 24.690 151.425 25.540 ;
        RECT 153.125 24.690 153.425 25.540 ;
        RECT 7.340 23.690 8.340 24.690 ;
        RECT 9.340 23.690 10.340 24.690 ;
        RECT 11.340 23.690 12.340 24.690 ;
        RECT 13.340 23.690 14.340 24.690 ;
        RECT 15.340 23.690 16.340 24.690 ;
        RECT 17.340 23.690 18.340 24.690 ;
        RECT 19.340 23.690 20.340 24.690 ;
        RECT 21.340 23.690 22.340 24.690 ;
        RECT 23.340 23.690 24.340 24.690 ;
        RECT 25.340 23.690 26.340 24.690 ;
        RECT 27.340 23.690 28.340 24.690 ;
        RECT 29.340 23.690 30.340 24.690 ;
        RECT 31.340 23.690 32.340 24.690 ;
        RECT 33.340 23.690 34.340 24.690 ;
        RECT 35.340 23.690 36.340 24.690 ;
        RECT 37.340 23.690 38.340 24.690 ;
        RECT 39.340 23.690 40.340 24.690 ;
        RECT 41.340 23.690 42.340 24.690 ;
        RECT 43.340 23.690 44.340 24.690 ;
        RECT 45.340 23.690 46.340 24.690 ;
        RECT 47.340 23.690 48.340 24.690 ;
        RECT 49.340 23.690 50.340 24.690 ;
        RECT 51.340 23.690 52.340 24.690 ;
        RECT 53.340 23.690 54.340 24.690 ;
        RECT 55.340 23.690 56.340 24.690 ;
        RECT 57.340 23.690 58.340 24.690 ;
        RECT 59.340 23.690 60.340 24.690 ;
        RECT 61.340 23.690 62.340 24.690 ;
        RECT 63.340 23.690 64.340 24.690 ;
        RECT 65.340 23.690 66.340 24.690 ;
        RECT 67.340 23.690 68.340 24.690 ;
        RECT 69.340 23.690 70.340 24.690 ;
        RECT 71.340 23.690 72.340 24.690 ;
        RECT 73.340 23.690 74.340 24.690 ;
        RECT 86.775 23.690 87.775 24.690 ;
        RECT 88.775 23.690 89.775 24.690 ;
        RECT 90.775 23.690 91.775 24.690 ;
        RECT 92.775 23.690 93.775 24.690 ;
        RECT 94.775 23.690 95.775 24.690 ;
        RECT 96.775 23.690 97.775 24.690 ;
        RECT 98.775 23.690 99.775 24.690 ;
        RECT 100.775 23.690 101.775 24.690 ;
        RECT 102.775 23.690 103.775 24.690 ;
        RECT 104.775 23.690 105.775 24.690 ;
        RECT 106.775 23.690 107.775 24.690 ;
        RECT 108.775 23.690 109.775 24.690 ;
        RECT 110.775 23.690 111.775 24.690 ;
        RECT 112.775 23.690 113.775 24.690 ;
        RECT 114.775 23.690 115.775 24.690 ;
        RECT 116.775 23.690 117.775 24.690 ;
        RECT 118.775 23.690 119.775 24.690 ;
        RECT 120.775 23.690 121.775 24.690 ;
        RECT 122.775 23.690 123.775 24.690 ;
        RECT 124.775 23.690 125.775 24.690 ;
        RECT 126.775 23.690 127.775 24.690 ;
        RECT 128.775 23.690 129.775 24.690 ;
        RECT 130.775 23.690 131.775 24.690 ;
        RECT 132.775 23.690 133.775 24.690 ;
        RECT 134.775 23.690 135.775 24.690 ;
        RECT 136.775 23.690 137.775 24.690 ;
        RECT 138.775 23.690 139.775 24.690 ;
        RECT 140.775 23.690 141.775 24.690 ;
        RECT 142.775 23.690 143.775 24.690 ;
        RECT 144.775 23.690 145.775 24.690 ;
        RECT 146.775 23.690 147.775 24.690 ;
        RECT 148.775 23.690 149.775 24.690 ;
        RECT 150.775 23.690 151.775 24.690 ;
        RECT 152.775 23.690 153.775 24.690 ;
        RECT 7.690 22.840 7.990 23.690 ;
        RECT 9.690 22.840 9.990 23.690 ;
        RECT 11.690 22.840 11.990 23.690 ;
        RECT 13.690 22.840 13.990 23.690 ;
        RECT 15.690 22.840 15.990 23.690 ;
        RECT 17.690 22.840 17.990 23.690 ;
        RECT 19.690 22.840 19.990 23.690 ;
        RECT 21.690 22.840 21.990 23.690 ;
        RECT 23.690 22.840 23.990 23.690 ;
        RECT 25.690 22.840 25.990 23.690 ;
        RECT 27.690 22.840 27.990 23.690 ;
        RECT 29.690 22.840 29.990 23.690 ;
        RECT 31.690 22.840 31.990 23.690 ;
        RECT 33.690 22.840 33.990 23.690 ;
        RECT 35.690 22.840 35.990 23.690 ;
        RECT 37.690 22.840 37.990 23.690 ;
        RECT 39.690 22.840 39.990 23.690 ;
        RECT 41.690 22.840 41.990 23.690 ;
        RECT 43.690 22.840 43.990 23.690 ;
        RECT 45.690 22.840 45.990 23.690 ;
        RECT 47.690 22.840 47.990 23.690 ;
        RECT 49.690 22.840 49.990 23.690 ;
        RECT 51.690 22.840 51.990 23.690 ;
        RECT 53.690 22.840 53.990 23.690 ;
        RECT 55.690 22.840 55.990 23.690 ;
        RECT 57.690 22.840 57.990 23.690 ;
        RECT 59.690 22.840 59.990 23.690 ;
        RECT 61.690 22.840 61.990 23.690 ;
        RECT 63.690 22.840 63.990 23.690 ;
        RECT 65.690 22.840 65.990 23.690 ;
        RECT 67.690 22.840 67.990 23.690 ;
        RECT 69.690 22.840 69.990 23.690 ;
        RECT 71.690 22.840 71.990 23.690 ;
        RECT 73.690 22.840 73.990 23.690 ;
        RECT 87.125 22.840 87.425 23.690 ;
        RECT 89.125 22.840 89.425 23.690 ;
        RECT 91.125 22.840 91.425 23.690 ;
        RECT 93.125 22.840 93.425 23.690 ;
        RECT 95.125 22.840 95.425 23.690 ;
        RECT 97.125 22.840 97.425 23.690 ;
        RECT 99.125 22.840 99.425 23.690 ;
        RECT 101.125 22.840 101.425 23.690 ;
        RECT 103.125 22.840 103.425 23.690 ;
        RECT 105.125 22.840 105.425 23.690 ;
        RECT 107.125 22.840 107.425 23.690 ;
        RECT 109.125 22.840 109.425 23.690 ;
        RECT 111.125 22.840 111.425 23.690 ;
        RECT 113.125 22.840 113.425 23.690 ;
        RECT 115.125 22.840 115.425 23.690 ;
        RECT 117.125 22.840 117.425 23.690 ;
        RECT 119.125 22.840 119.425 23.690 ;
        RECT 121.125 22.840 121.425 23.690 ;
        RECT 123.125 22.840 123.425 23.690 ;
        RECT 125.125 22.840 125.425 23.690 ;
        RECT 127.125 22.840 127.425 23.690 ;
        RECT 129.125 22.840 129.425 23.690 ;
        RECT 131.125 22.840 131.425 23.690 ;
        RECT 133.125 22.840 133.425 23.690 ;
        RECT 135.125 22.840 135.425 23.690 ;
        RECT 137.125 22.840 137.425 23.690 ;
        RECT 139.125 22.840 139.425 23.690 ;
        RECT 141.125 22.840 141.425 23.690 ;
        RECT 143.125 22.840 143.425 23.690 ;
        RECT 145.125 22.840 145.425 23.690 ;
        RECT 147.125 22.840 147.425 23.690 ;
        RECT 149.125 22.840 149.425 23.690 ;
        RECT 151.125 22.840 151.425 23.690 ;
        RECT 153.125 22.840 153.425 23.690 ;
        RECT 7.340 21.840 8.340 22.840 ;
        RECT 9.340 21.840 10.340 22.840 ;
        RECT 11.340 21.840 12.340 22.840 ;
        RECT 13.340 21.840 14.340 22.840 ;
        RECT 15.340 21.840 16.340 22.840 ;
        RECT 17.340 21.840 18.340 22.840 ;
        RECT 19.340 21.840 20.340 22.840 ;
        RECT 21.340 21.840 22.340 22.840 ;
        RECT 23.340 21.840 24.340 22.840 ;
        RECT 25.340 21.840 26.340 22.840 ;
        RECT 27.340 21.840 28.340 22.840 ;
        RECT 29.340 21.840 30.340 22.840 ;
        RECT 31.340 21.840 32.340 22.840 ;
        RECT 33.340 21.840 34.340 22.840 ;
        RECT 35.340 21.840 36.340 22.840 ;
        RECT 37.340 21.840 38.340 22.840 ;
        RECT 39.340 21.840 40.340 22.840 ;
        RECT 41.340 21.840 42.340 22.840 ;
        RECT 43.340 21.840 44.340 22.840 ;
        RECT 45.340 21.840 46.340 22.840 ;
        RECT 47.340 21.840 48.340 22.840 ;
        RECT 49.340 21.840 50.340 22.840 ;
        RECT 51.340 21.840 52.340 22.840 ;
        RECT 53.340 21.840 54.340 22.840 ;
        RECT 55.340 21.840 56.340 22.840 ;
        RECT 57.340 21.840 58.340 22.840 ;
        RECT 59.340 21.840 60.340 22.840 ;
        RECT 61.340 21.840 62.340 22.840 ;
        RECT 63.340 21.840 64.340 22.840 ;
        RECT 65.340 21.840 66.340 22.840 ;
        RECT 67.340 21.840 68.340 22.840 ;
        RECT 69.340 21.840 70.340 22.840 ;
        RECT 71.340 21.840 72.340 22.840 ;
        RECT 73.340 21.840 74.340 22.840 ;
        RECT 86.775 21.840 87.775 22.840 ;
        RECT 88.775 21.840 89.775 22.840 ;
        RECT 90.775 21.840 91.775 22.840 ;
        RECT 92.775 21.840 93.775 22.840 ;
        RECT 94.775 21.840 95.775 22.840 ;
        RECT 96.775 21.840 97.775 22.840 ;
        RECT 98.775 21.840 99.775 22.840 ;
        RECT 100.775 21.840 101.775 22.840 ;
        RECT 102.775 21.840 103.775 22.840 ;
        RECT 104.775 21.840 105.775 22.840 ;
        RECT 106.775 21.840 107.775 22.840 ;
        RECT 108.775 21.840 109.775 22.840 ;
        RECT 110.775 21.840 111.775 22.840 ;
        RECT 112.775 21.840 113.775 22.840 ;
        RECT 114.775 21.840 115.775 22.840 ;
        RECT 116.775 21.840 117.775 22.840 ;
        RECT 118.775 21.840 119.775 22.840 ;
        RECT 120.775 21.840 121.775 22.840 ;
        RECT 122.775 21.840 123.775 22.840 ;
        RECT 124.775 21.840 125.775 22.840 ;
        RECT 126.775 21.840 127.775 22.840 ;
        RECT 128.775 21.840 129.775 22.840 ;
        RECT 130.775 21.840 131.775 22.840 ;
        RECT 132.775 21.840 133.775 22.840 ;
        RECT 134.775 21.840 135.775 22.840 ;
        RECT 136.775 21.840 137.775 22.840 ;
        RECT 138.775 21.840 139.775 22.840 ;
        RECT 140.775 21.840 141.775 22.840 ;
        RECT 142.775 21.840 143.775 22.840 ;
        RECT 144.775 21.840 145.775 22.840 ;
        RECT 146.775 21.840 147.775 22.840 ;
        RECT 148.775 21.840 149.775 22.840 ;
        RECT 150.775 21.840 151.775 22.840 ;
        RECT 152.775 21.840 153.775 22.840 ;
        RECT 7.690 20.990 7.990 21.840 ;
        RECT 9.690 20.990 9.990 21.840 ;
        RECT 11.690 20.990 11.990 21.840 ;
        RECT 13.690 20.990 13.990 21.840 ;
        RECT 15.690 20.990 15.990 21.840 ;
        RECT 17.690 20.990 17.990 21.840 ;
        RECT 19.690 20.990 19.990 21.840 ;
        RECT 21.690 20.990 21.990 21.840 ;
        RECT 23.690 20.990 23.990 21.840 ;
        RECT 25.690 20.990 25.990 21.840 ;
        RECT 27.690 20.990 27.990 21.840 ;
        RECT 29.690 20.990 29.990 21.840 ;
        RECT 31.690 20.990 31.990 21.840 ;
        RECT 33.690 20.990 33.990 21.840 ;
        RECT 35.690 20.990 35.990 21.840 ;
        RECT 37.690 20.990 37.990 21.840 ;
        RECT 39.690 20.990 39.990 21.840 ;
        RECT 41.690 20.990 41.990 21.840 ;
        RECT 43.690 20.990 43.990 21.840 ;
        RECT 45.690 20.990 45.990 21.840 ;
        RECT 47.690 20.990 47.990 21.840 ;
        RECT 49.690 20.990 49.990 21.840 ;
        RECT 51.690 20.990 51.990 21.840 ;
        RECT 53.690 20.990 53.990 21.840 ;
        RECT 55.690 20.990 55.990 21.840 ;
        RECT 57.690 20.990 57.990 21.840 ;
        RECT 59.690 20.990 59.990 21.840 ;
        RECT 61.690 20.990 61.990 21.840 ;
        RECT 63.690 20.990 63.990 21.840 ;
        RECT 65.690 20.990 65.990 21.840 ;
        RECT 67.690 20.990 67.990 21.840 ;
        RECT 69.690 20.990 69.990 21.840 ;
        RECT 71.690 20.990 71.990 21.840 ;
        RECT 73.690 20.990 73.990 21.840 ;
        RECT 87.125 20.990 87.425 21.840 ;
        RECT 89.125 20.990 89.425 21.840 ;
        RECT 91.125 20.990 91.425 21.840 ;
        RECT 93.125 20.990 93.425 21.840 ;
        RECT 95.125 20.990 95.425 21.840 ;
        RECT 97.125 20.990 97.425 21.840 ;
        RECT 99.125 20.990 99.425 21.840 ;
        RECT 101.125 20.990 101.425 21.840 ;
        RECT 103.125 20.990 103.425 21.840 ;
        RECT 105.125 20.990 105.425 21.840 ;
        RECT 107.125 20.990 107.425 21.840 ;
        RECT 109.125 20.990 109.425 21.840 ;
        RECT 111.125 20.990 111.425 21.840 ;
        RECT 113.125 20.990 113.425 21.840 ;
        RECT 115.125 20.990 115.425 21.840 ;
        RECT 117.125 20.990 117.425 21.840 ;
        RECT 119.125 20.990 119.425 21.840 ;
        RECT 121.125 20.990 121.425 21.840 ;
        RECT 123.125 20.990 123.425 21.840 ;
        RECT 125.125 20.990 125.425 21.840 ;
        RECT 127.125 20.990 127.425 21.840 ;
        RECT 129.125 20.990 129.425 21.840 ;
        RECT 131.125 20.990 131.425 21.840 ;
        RECT 133.125 20.990 133.425 21.840 ;
        RECT 135.125 20.990 135.425 21.840 ;
        RECT 137.125 20.990 137.425 21.840 ;
        RECT 139.125 20.990 139.425 21.840 ;
        RECT 141.125 20.990 141.425 21.840 ;
        RECT 143.125 20.990 143.425 21.840 ;
        RECT 145.125 20.990 145.425 21.840 ;
        RECT 147.125 20.990 147.425 21.840 ;
        RECT 149.125 20.990 149.425 21.840 ;
        RECT 151.125 20.990 151.425 21.840 ;
        RECT 153.125 20.990 153.425 21.840 ;
        RECT 7.340 19.990 8.340 20.990 ;
        RECT 9.340 19.990 10.340 20.990 ;
        RECT 11.340 19.990 12.340 20.990 ;
        RECT 13.340 19.990 14.340 20.990 ;
        RECT 15.340 19.990 16.340 20.990 ;
        RECT 17.340 19.990 18.340 20.990 ;
        RECT 19.340 19.990 20.340 20.990 ;
        RECT 21.340 19.990 22.340 20.990 ;
        RECT 23.340 19.990 24.340 20.990 ;
        RECT 25.340 19.990 26.340 20.990 ;
        RECT 27.340 19.990 28.340 20.990 ;
        RECT 29.340 19.990 30.340 20.990 ;
        RECT 31.340 19.990 32.340 20.990 ;
        RECT 33.340 19.990 34.340 20.990 ;
        RECT 35.340 19.990 36.340 20.990 ;
        RECT 37.340 19.990 38.340 20.990 ;
        RECT 39.340 19.990 40.340 20.990 ;
        RECT 41.340 19.990 42.340 20.990 ;
        RECT 43.340 19.990 44.340 20.990 ;
        RECT 45.340 19.990 46.340 20.990 ;
        RECT 47.340 19.990 48.340 20.990 ;
        RECT 49.340 19.990 50.340 20.990 ;
        RECT 51.340 19.990 52.340 20.990 ;
        RECT 53.340 19.990 54.340 20.990 ;
        RECT 55.340 19.990 56.340 20.990 ;
        RECT 57.340 19.990 58.340 20.990 ;
        RECT 59.340 19.990 60.340 20.990 ;
        RECT 61.340 19.990 62.340 20.990 ;
        RECT 63.340 19.990 64.340 20.990 ;
        RECT 65.340 19.990 66.340 20.990 ;
        RECT 67.340 19.990 68.340 20.990 ;
        RECT 69.340 19.990 70.340 20.990 ;
        RECT 71.340 19.990 72.340 20.990 ;
        RECT 73.340 19.990 74.340 20.990 ;
        RECT 86.775 19.990 87.775 20.990 ;
        RECT 88.775 19.990 89.775 20.990 ;
        RECT 90.775 19.990 91.775 20.990 ;
        RECT 92.775 19.990 93.775 20.990 ;
        RECT 94.775 19.990 95.775 20.990 ;
        RECT 96.775 19.990 97.775 20.990 ;
        RECT 98.775 19.990 99.775 20.990 ;
        RECT 100.775 19.990 101.775 20.990 ;
        RECT 102.775 19.990 103.775 20.990 ;
        RECT 104.775 19.990 105.775 20.990 ;
        RECT 106.775 19.990 107.775 20.990 ;
        RECT 108.775 19.990 109.775 20.990 ;
        RECT 110.775 19.990 111.775 20.990 ;
        RECT 112.775 19.990 113.775 20.990 ;
        RECT 114.775 19.990 115.775 20.990 ;
        RECT 116.775 19.990 117.775 20.990 ;
        RECT 118.775 19.990 119.775 20.990 ;
        RECT 120.775 19.990 121.775 20.990 ;
        RECT 122.775 19.990 123.775 20.990 ;
        RECT 124.775 19.990 125.775 20.990 ;
        RECT 126.775 19.990 127.775 20.990 ;
        RECT 128.775 19.990 129.775 20.990 ;
        RECT 130.775 19.990 131.775 20.990 ;
        RECT 132.775 19.990 133.775 20.990 ;
        RECT 134.775 19.990 135.775 20.990 ;
        RECT 136.775 19.990 137.775 20.990 ;
        RECT 138.775 19.990 139.775 20.990 ;
        RECT 140.775 19.990 141.775 20.990 ;
        RECT 142.775 19.990 143.775 20.990 ;
        RECT 144.775 19.990 145.775 20.990 ;
        RECT 146.775 19.990 147.775 20.990 ;
        RECT 148.775 19.990 149.775 20.990 ;
        RECT 150.775 19.990 151.775 20.990 ;
        RECT 152.775 19.990 153.775 20.990 ;
        RECT 7.690 19.140 7.990 19.990 ;
        RECT 9.690 19.140 9.990 19.990 ;
        RECT 11.690 19.140 11.990 19.990 ;
        RECT 13.690 19.140 13.990 19.990 ;
        RECT 15.690 19.140 15.990 19.990 ;
        RECT 17.690 19.140 17.990 19.990 ;
        RECT 19.690 19.140 19.990 19.990 ;
        RECT 21.690 19.140 21.990 19.990 ;
        RECT 23.690 19.140 23.990 19.990 ;
        RECT 25.690 19.140 25.990 19.990 ;
        RECT 27.690 19.140 27.990 19.990 ;
        RECT 29.690 19.140 29.990 19.990 ;
        RECT 31.690 19.140 31.990 19.990 ;
        RECT 33.690 19.140 33.990 19.990 ;
        RECT 35.690 19.140 35.990 19.990 ;
        RECT 37.690 19.140 37.990 19.990 ;
        RECT 39.690 19.140 39.990 19.990 ;
        RECT 41.690 19.140 41.990 19.990 ;
        RECT 43.690 19.140 43.990 19.990 ;
        RECT 45.690 19.140 45.990 19.990 ;
        RECT 47.690 19.140 47.990 19.990 ;
        RECT 49.690 19.140 49.990 19.990 ;
        RECT 51.690 19.140 51.990 19.990 ;
        RECT 53.690 19.140 53.990 19.990 ;
        RECT 55.690 19.140 55.990 19.990 ;
        RECT 57.690 19.140 57.990 19.990 ;
        RECT 59.690 19.140 59.990 19.990 ;
        RECT 61.690 19.140 61.990 19.990 ;
        RECT 63.690 19.140 63.990 19.990 ;
        RECT 65.690 19.140 65.990 19.990 ;
        RECT 67.690 19.140 67.990 19.990 ;
        RECT 69.690 19.140 69.990 19.990 ;
        RECT 71.690 19.140 71.990 19.990 ;
        RECT 73.690 19.140 73.990 19.990 ;
        RECT 87.125 19.140 87.425 19.990 ;
        RECT 89.125 19.140 89.425 19.990 ;
        RECT 91.125 19.140 91.425 19.990 ;
        RECT 93.125 19.140 93.425 19.990 ;
        RECT 95.125 19.140 95.425 19.990 ;
        RECT 97.125 19.140 97.425 19.990 ;
        RECT 99.125 19.140 99.425 19.990 ;
        RECT 101.125 19.140 101.425 19.990 ;
        RECT 103.125 19.140 103.425 19.990 ;
        RECT 105.125 19.140 105.425 19.990 ;
        RECT 107.125 19.140 107.425 19.990 ;
        RECT 109.125 19.140 109.425 19.990 ;
        RECT 111.125 19.140 111.425 19.990 ;
        RECT 113.125 19.140 113.425 19.990 ;
        RECT 115.125 19.140 115.425 19.990 ;
        RECT 117.125 19.140 117.425 19.990 ;
        RECT 119.125 19.140 119.425 19.990 ;
        RECT 121.125 19.140 121.425 19.990 ;
        RECT 123.125 19.140 123.425 19.990 ;
        RECT 125.125 19.140 125.425 19.990 ;
        RECT 127.125 19.140 127.425 19.990 ;
        RECT 129.125 19.140 129.425 19.990 ;
        RECT 131.125 19.140 131.425 19.990 ;
        RECT 133.125 19.140 133.425 19.990 ;
        RECT 135.125 19.140 135.425 19.990 ;
        RECT 137.125 19.140 137.425 19.990 ;
        RECT 139.125 19.140 139.425 19.990 ;
        RECT 141.125 19.140 141.425 19.990 ;
        RECT 143.125 19.140 143.425 19.990 ;
        RECT 145.125 19.140 145.425 19.990 ;
        RECT 147.125 19.140 147.425 19.990 ;
        RECT 149.125 19.140 149.425 19.990 ;
        RECT 151.125 19.140 151.425 19.990 ;
        RECT 153.125 19.140 153.425 19.990 ;
        RECT 7.340 18.140 8.340 19.140 ;
        RECT 9.340 18.140 10.340 19.140 ;
        RECT 11.340 18.140 12.340 19.140 ;
        RECT 13.340 18.140 14.340 19.140 ;
        RECT 15.340 18.140 16.340 19.140 ;
        RECT 17.340 18.140 18.340 19.140 ;
        RECT 19.340 18.140 20.340 19.140 ;
        RECT 21.340 18.140 22.340 19.140 ;
        RECT 23.340 18.140 24.340 19.140 ;
        RECT 25.340 18.140 26.340 19.140 ;
        RECT 27.340 18.140 28.340 19.140 ;
        RECT 29.340 18.140 30.340 19.140 ;
        RECT 31.340 18.140 32.340 19.140 ;
        RECT 33.340 18.140 34.340 19.140 ;
        RECT 35.340 18.140 36.340 19.140 ;
        RECT 37.340 18.140 38.340 19.140 ;
        RECT 39.340 18.140 40.340 19.140 ;
        RECT 41.340 18.140 42.340 19.140 ;
        RECT 43.340 18.140 44.340 19.140 ;
        RECT 45.340 18.140 46.340 19.140 ;
        RECT 47.340 18.140 48.340 19.140 ;
        RECT 49.340 18.140 50.340 19.140 ;
        RECT 51.340 18.140 52.340 19.140 ;
        RECT 53.340 18.140 54.340 19.140 ;
        RECT 55.340 18.140 56.340 19.140 ;
        RECT 57.340 18.140 58.340 19.140 ;
        RECT 59.340 18.140 60.340 19.140 ;
        RECT 61.340 18.140 62.340 19.140 ;
        RECT 63.340 18.140 64.340 19.140 ;
        RECT 65.340 18.140 66.340 19.140 ;
        RECT 67.340 18.140 68.340 19.140 ;
        RECT 69.340 18.140 70.340 19.140 ;
        RECT 71.340 18.140 72.340 19.140 ;
        RECT 73.340 18.140 74.340 19.140 ;
        RECT 86.775 18.140 87.775 19.140 ;
        RECT 88.775 18.140 89.775 19.140 ;
        RECT 90.775 18.140 91.775 19.140 ;
        RECT 92.775 18.140 93.775 19.140 ;
        RECT 94.775 18.140 95.775 19.140 ;
        RECT 96.775 18.140 97.775 19.140 ;
        RECT 98.775 18.140 99.775 19.140 ;
        RECT 100.775 18.140 101.775 19.140 ;
        RECT 102.775 18.140 103.775 19.140 ;
        RECT 104.775 18.140 105.775 19.140 ;
        RECT 106.775 18.140 107.775 19.140 ;
        RECT 108.775 18.140 109.775 19.140 ;
        RECT 110.775 18.140 111.775 19.140 ;
        RECT 112.775 18.140 113.775 19.140 ;
        RECT 114.775 18.140 115.775 19.140 ;
        RECT 116.775 18.140 117.775 19.140 ;
        RECT 118.775 18.140 119.775 19.140 ;
        RECT 120.775 18.140 121.775 19.140 ;
        RECT 122.775 18.140 123.775 19.140 ;
        RECT 124.775 18.140 125.775 19.140 ;
        RECT 126.775 18.140 127.775 19.140 ;
        RECT 128.775 18.140 129.775 19.140 ;
        RECT 130.775 18.140 131.775 19.140 ;
        RECT 132.775 18.140 133.775 19.140 ;
        RECT 134.775 18.140 135.775 19.140 ;
        RECT 136.775 18.140 137.775 19.140 ;
        RECT 138.775 18.140 139.775 19.140 ;
        RECT 140.775 18.140 141.775 19.140 ;
        RECT 142.775 18.140 143.775 19.140 ;
        RECT 144.775 18.140 145.775 19.140 ;
        RECT 146.775 18.140 147.775 19.140 ;
        RECT 148.775 18.140 149.775 19.140 ;
        RECT 150.775 18.140 151.775 19.140 ;
        RECT 152.775 18.140 153.775 19.140 ;
        RECT 7.690 17.290 7.990 18.140 ;
        RECT 9.690 17.290 9.990 18.140 ;
        RECT 11.690 17.290 11.990 18.140 ;
        RECT 13.690 17.290 13.990 18.140 ;
        RECT 15.690 17.290 15.990 18.140 ;
        RECT 17.690 17.290 17.990 18.140 ;
        RECT 19.690 17.290 19.990 18.140 ;
        RECT 21.690 17.290 21.990 18.140 ;
        RECT 23.690 17.290 23.990 18.140 ;
        RECT 25.690 17.290 25.990 18.140 ;
        RECT 27.690 17.290 27.990 18.140 ;
        RECT 29.690 17.290 29.990 18.140 ;
        RECT 31.690 17.290 31.990 18.140 ;
        RECT 33.690 17.290 33.990 18.140 ;
        RECT 35.690 17.290 35.990 18.140 ;
        RECT 37.690 17.290 37.990 18.140 ;
        RECT 39.690 17.290 39.990 18.140 ;
        RECT 41.690 17.290 41.990 18.140 ;
        RECT 43.690 17.290 43.990 18.140 ;
        RECT 45.690 17.290 45.990 18.140 ;
        RECT 47.690 17.290 47.990 18.140 ;
        RECT 49.690 17.290 49.990 18.140 ;
        RECT 51.690 17.290 51.990 18.140 ;
        RECT 53.690 17.290 53.990 18.140 ;
        RECT 55.690 17.290 55.990 18.140 ;
        RECT 57.690 17.290 57.990 18.140 ;
        RECT 59.690 17.290 59.990 18.140 ;
        RECT 61.690 17.290 61.990 18.140 ;
        RECT 63.690 17.290 63.990 18.140 ;
        RECT 65.690 17.290 65.990 18.140 ;
        RECT 67.690 17.290 67.990 18.140 ;
        RECT 69.690 17.290 69.990 18.140 ;
        RECT 71.690 17.290 71.990 18.140 ;
        RECT 73.690 17.290 73.990 18.140 ;
        RECT 87.125 17.290 87.425 18.140 ;
        RECT 89.125 17.290 89.425 18.140 ;
        RECT 91.125 17.290 91.425 18.140 ;
        RECT 93.125 17.290 93.425 18.140 ;
        RECT 95.125 17.290 95.425 18.140 ;
        RECT 97.125 17.290 97.425 18.140 ;
        RECT 99.125 17.290 99.425 18.140 ;
        RECT 101.125 17.290 101.425 18.140 ;
        RECT 103.125 17.290 103.425 18.140 ;
        RECT 105.125 17.290 105.425 18.140 ;
        RECT 107.125 17.290 107.425 18.140 ;
        RECT 109.125 17.290 109.425 18.140 ;
        RECT 111.125 17.290 111.425 18.140 ;
        RECT 113.125 17.290 113.425 18.140 ;
        RECT 115.125 17.290 115.425 18.140 ;
        RECT 117.125 17.290 117.425 18.140 ;
        RECT 119.125 17.290 119.425 18.140 ;
        RECT 121.125 17.290 121.425 18.140 ;
        RECT 123.125 17.290 123.425 18.140 ;
        RECT 125.125 17.290 125.425 18.140 ;
        RECT 127.125 17.290 127.425 18.140 ;
        RECT 129.125 17.290 129.425 18.140 ;
        RECT 131.125 17.290 131.425 18.140 ;
        RECT 133.125 17.290 133.425 18.140 ;
        RECT 135.125 17.290 135.425 18.140 ;
        RECT 137.125 17.290 137.425 18.140 ;
        RECT 139.125 17.290 139.425 18.140 ;
        RECT 141.125 17.290 141.425 18.140 ;
        RECT 143.125 17.290 143.425 18.140 ;
        RECT 145.125 17.290 145.425 18.140 ;
        RECT 147.125 17.290 147.425 18.140 ;
        RECT 149.125 17.290 149.425 18.140 ;
        RECT 151.125 17.290 151.425 18.140 ;
        RECT 153.125 17.290 153.425 18.140 ;
        RECT 7.340 16.290 8.340 17.290 ;
        RECT 9.340 16.290 10.340 17.290 ;
        RECT 11.340 16.290 12.340 17.290 ;
        RECT 13.340 16.290 14.340 17.290 ;
        RECT 15.340 16.290 16.340 17.290 ;
        RECT 17.340 16.290 18.340 17.290 ;
        RECT 19.340 16.290 20.340 17.290 ;
        RECT 21.340 16.290 22.340 17.290 ;
        RECT 23.340 16.290 24.340 17.290 ;
        RECT 25.340 16.290 26.340 17.290 ;
        RECT 27.340 16.290 28.340 17.290 ;
        RECT 29.340 16.290 30.340 17.290 ;
        RECT 31.340 16.290 32.340 17.290 ;
        RECT 33.340 16.290 34.340 17.290 ;
        RECT 35.340 16.290 36.340 17.290 ;
        RECT 37.340 16.290 38.340 17.290 ;
        RECT 39.340 16.290 40.340 17.290 ;
        RECT 41.340 16.290 42.340 17.290 ;
        RECT 43.340 16.290 44.340 17.290 ;
        RECT 45.340 16.290 46.340 17.290 ;
        RECT 47.340 16.290 48.340 17.290 ;
        RECT 49.340 16.290 50.340 17.290 ;
        RECT 51.340 16.290 52.340 17.290 ;
        RECT 53.340 16.290 54.340 17.290 ;
        RECT 55.340 16.290 56.340 17.290 ;
        RECT 57.340 16.290 58.340 17.290 ;
        RECT 59.340 16.290 60.340 17.290 ;
        RECT 61.340 16.290 62.340 17.290 ;
        RECT 63.340 16.290 64.340 17.290 ;
        RECT 65.340 16.290 66.340 17.290 ;
        RECT 67.340 16.290 68.340 17.290 ;
        RECT 69.340 16.290 70.340 17.290 ;
        RECT 71.340 16.290 72.340 17.290 ;
        RECT 73.340 16.290 74.340 17.290 ;
        RECT 86.775 16.290 87.775 17.290 ;
        RECT 88.775 16.290 89.775 17.290 ;
        RECT 90.775 16.290 91.775 17.290 ;
        RECT 92.775 16.290 93.775 17.290 ;
        RECT 94.775 16.290 95.775 17.290 ;
        RECT 96.775 16.290 97.775 17.290 ;
        RECT 98.775 16.290 99.775 17.290 ;
        RECT 100.775 16.290 101.775 17.290 ;
        RECT 102.775 16.290 103.775 17.290 ;
        RECT 104.775 16.290 105.775 17.290 ;
        RECT 106.775 16.290 107.775 17.290 ;
        RECT 108.775 16.290 109.775 17.290 ;
        RECT 110.775 16.290 111.775 17.290 ;
        RECT 112.775 16.290 113.775 17.290 ;
        RECT 114.775 16.290 115.775 17.290 ;
        RECT 116.775 16.290 117.775 17.290 ;
        RECT 118.775 16.290 119.775 17.290 ;
        RECT 120.775 16.290 121.775 17.290 ;
        RECT 122.775 16.290 123.775 17.290 ;
        RECT 124.775 16.290 125.775 17.290 ;
        RECT 126.775 16.290 127.775 17.290 ;
        RECT 128.775 16.290 129.775 17.290 ;
        RECT 130.775 16.290 131.775 17.290 ;
        RECT 132.775 16.290 133.775 17.290 ;
        RECT 134.775 16.290 135.775 17.290 ;
        RECT 136.775 16.290 137.775 17.290 ;
        RECT 138.775 16.290 139.775 17.290 ;
        RECT 140.775 16.290 141.775 17.290 ;
        RECT 142.775 16.290 143.775 17.290 ;
        RECT 144.775 16.290 145.775 17.290 ;
        RECT 146.775 16.290 147.775 17.290 ;
        RECT 148.775 16.290 149.775 17.290 ;
        RECT 150.775 16.290 151.775 17.290 ;
        RECT 152.775 16.290 153.775 17.290 ;
        RECT 7.690 15.440 7.990 16.290 ;
        RECT 9.690 15.440 9.990 16.290 ;
        RECT 11.690 15.440 11.990 16.290 ;
        RECT 13.690 15.440 13.990 16.290 ;
        RECT 15.690 15.440 15.990 16.290 ;
        RECT 17.690 15.440 17.990 16.290 ;
        RECT 19.690 15.440 19.990 16.290 ;
        RECT 21.690 15.440 21.990 16.290 ;
        RECT 23.690 15.440 23.990 16.290 ;
        RECT 25.690 15.440 25.990 16.290 ;
        RECT 27.690 15.440 27.990 16.290 ;
        RECT 29.690 15.440 29.990 16.290 ;
        RECT 31.690 15.440 31.990 16.290 ;
        RECT 33.690 15.440 33.990 16.290 ;
        RECT 35.690 15.440 35.990 16.290 ;
        RECT 37.690 15.440 37.990 16.290 ;
        RECT 39.690 15.440 39.990 16.290 ;
        RECT 41.690 15.440 41.990 16.290 ;
        RECT 43.690 15.440 43.990 16.290 ;
        RECT 45.690 15.440 45.990 16.290 ;
        RECT 47.690 15.440 47.990 16.290 ;
        RECT 49.690 15.440 49.990 16.290 ;
        RECT 51.690 15.440 51.990 16.290 ;
        RECT 53.690 15.440 53.990 16.290 ;
        RECT 55.690 15.440 55.990 16.290 ;
        RECT 57.690 15.440 57.990 16.290 ;
        RECT 59.690 15.440 59.990 16.290 ;
        RECT 61.690 15.440 61.990 16.290 ;
        RECT 63.690 15.440 63.990 16.290 ;
        RECT 65.690 15.440 65.990 16.290 ;
        RECT 67.690 15.440 67.990 16.290 ;
        RECT 69.690 15.440 69.990 16.290 ;
        RECT 71.690 15.440 71.990 16.290 ;
        RECT 73.690 15.440 73.990 16.290 ;
        RECT 87.125 15.440 87.425 16.290 ;
        RECT 89.125 15.440 89.425 16.290 ;
        RECT 91.125 15.440 91.425 16.290 ;
        RECT 93.125 15.440 93.425 16.290 ;
        RECT 95.125 15.440 95.425 16.290 ;
        RECT 97.125 15.440 97.425 16.290 ;
        RECT 99.125 15.440 99.425 16.290 ;
        RECT 101.125 15.440 101.425 16.290 ;
        RECT 103.125 15.440 103.425 16.290 ;
        RECT 105.125 15.440 105.425 16.290 ;
        RECT 107.125 15.440 107.425 16.290 ;
        RECT 109.125 15.440 109.425 16.290 ;
        RECT 111.125 15.440 111.425 16.290 ;
        RECT 113.125 15.440 113.425 16.290 ;
        RECT 115.125 15.440 115.425 16.290 ;
        RECT 117.125 15.440 117.425 16.290 ;
        RECT 119.125 15.440 119.425 16.290 ;
        RECT 121.125 15.440 121.425 16.290 ;
        RECT 123.125 15.440 123.425 16.290 ;
        RECT 125.125 15.440 125.425 16.290 ;
        RECT 127.125 15.440 127.425 16.290 ;
        RECT 129.125 15.440 129.425 16.290 ;
        RECT 131.125 15.440 131.425 16.290 ;
        RECT 133.125 15.440 133.425 16.290 ;
        RECT 135.125 15.440 135.425 16.290 ;
        RECT 137.125 15.440 137.425 16.290 ;
        RECT 139.125 15.440 139.425 16.290 ;
        RECT 141.125 15.440 141.425 16.290 ;
        RECT 143.125 15.440 143.425 16.290 ;
        RECT 145.125 15.440 145.425 16.290 ;
        RECT 147.125 15.440 147.425 16.290 ;
        RECT 149.125 15.440 149.425 16.290 ;
        RECT 151.125 15.440 151.425 16.290 ;
        RECT 153.125 15.440 153.425 16.290 ;
        RECT 7.340 14.440 8.340 15.440 ;
        RECT 9.340 14.440 10.340 15.440 ;
        RECT 11.340 14.440 12.340 15.440 ;
        RECT 13.340 14.440 14.340 15.440 ;
        RECT 15.340 14.440 16.340 15.440 ;
        RECT 17.340 14.440 18.340 15.440 ;
        RECT 19.340 14.440 20.340 15.440 ;
        RECT 21.340 14.440 22.340 15.440 ;
        RECT 23.340 14.440 24.340 15.440 ;
        RECT 25.340 14.440 26.340 15.440 ;
        RECT 27.340 14.440 28.340 15.440 ;
        RECT 29.340 14.440 30.340 15.440 ;
        RECT 31.340 14.440 32.340 15.440 ;
        RECT 33.340 14.440 34.340 15.440 ;
        RECT 35.340 14.440 36.340 15.440 ;
        RECT 37.340 14.440 38.340 15.440 ;
        RECT 39.340 14.440 40.340 15.440 ;
        RECT 41.340 14.440 42.340 15.440 ;
        RECT 43.340 14.440 44.340 15.440 ;
        RECT 45.340 14.440 46.340 15.440 ;
        RECT 47.340 14.440 48.340 15.440 ;
        RECT 49.340 14.440 50.340 15.440 ;
        RECT 51.340 14.440 52.340 15.440 ;
        RECT 53.340 14.440 54.340 15.440 ;
        RECT 55.340 14.440 56.340 15.440 ;
        RECT 57.340 14.440 58.340 15.440 ;
        RECT 59.340 14.440 60.340 15.440 ;
        RECT 61.340 14.440 62.340 15.440 ;
        RECT 63.340 14.440 64.340 15.440 ;
        RECT 65.340 14.440 66.340 15.440 ;
        RECT 67.340 14.440 68.340 15.440 ;
        RECT 69.340 14.440 70.340 15.440 ;
        RECT 71.340 14.440 72.340 15.440 ;
        RECT 73.340 14.440 74.340 15.440 ;
        RECT 86.775 14.440 87.775 15.440 ;
        RECT 88.775 14.440 89.775 15.440 ;
        RECT 90.775 14.440 91.775 15.440 ;
        RECT 92.775 14.440 93.775 15.440 ;
        RECT 94.775 14.440 95.775 15.440 ;
        RECT 96.775 14.440 97.775 15.440 ;
        RECT 98.775 14.440 99.775 15.440 ;
        RECT 100.775 14.440 101.775 15.440 ;
        RECT 102.775 14.440 103.775 15.440 ;
        RECT 104.775 14.440 105.775 15.440 ;
        RECT 106.775 14.440 107.775 15.440 ;
        RECT 108.775 14.440 109.775 15.440 ;
        RECT 110.775 14.440 111.775 15.440 ;
        RECT 112.775 14.440 113.775 15.440 ;
        RECT 114.775 14.440 115.775 15.440 ;
        RECT 116.775 14.440 117.775 15.440 ;
        RECT 118.775 14.440 119.775 15.440 ;
        RECT 120.775 14.440 121.775 15.440 ;
        RECT 122.775 14.440 123.775 15.440 ;
        RECT 124.775 14.440 125.775 15.440 ;
        RECT 126.775 14.440 127.775 15.440 ;
        RECT 128.775 14.440 129.775 15.440 ;
        RECT 130.775 14.440 131.775 15.440 ;
        RECT 132.775 14.440 133.775 15.440 ;
        RECT 134.775 14.440 135.775 15.440 ;
        RECT 136.775 14.440 137.775 15.440 ;
        RECT 138.775 14.440 139.775 15.440 ;
        RECT 140.775 14.440 141.775 15.440 ;
        RECT 142.775 14.440 143.775 15.440 ;
        RECT 144.775 14.440 145.775 15.440 ;
        RECT 146.775 14.440 147.775 15.440 ;
        RECT 148.775 14.440 149.775 15.440 ;
        RECT 150.775 14.440 151.775 15.440 ;
        RECT 152.775 14.440 153.775 15.440 ;
        RECT 7.690 13.590 7.990 14.440 ;
        RECT 9.690 13.590 9.990 14.440 ;
        RECT 11.690 13.590 11.990 14.440 ;
        RECT 13.690 13.590 13.990 14.440 ;
        RECT 15.690 13.590 15.990 14.440 ;
        RECT 17.690 13.590 17.990 14.440 ;
        RECT 19.690 13.590 19.990 14.440 ;
        RECT 21.690 13.590 21.990 14.440 ;
        RECT 23.690 13.590 23.990 14.440 ;
        RECT 25.690 13.590 25.990 14.440 ;
        RECT 27.690 13.590 27.990 14.440 ;
        RECT 29.690 13.590 29.990 14.440 ;
        RECT 31.690 13.590 31.990 14.440 ;
        RECT 33.690 13.590 33.990 14.440 ;
        RECT 35.690 13.590 35.990 14.440 ;
        RECT 37.690 13.590 37.990 14.440 ;
        RECT 39.690 13.590 39.990 14.440 ;
        RECT 41.690 13.590 41.990 14.440 ;
        RECT 43.690 13.590 43.990 14.440 ;
        RECT 45.690 13.590 45.990 14.440 ;
        RECT 47.690 13.590 47.990 14.440 ;
        RECT 49.690 13.590 49.990 14.440 ;
        RECT 51.690 13.590 51.990 14.440 ;
        RECT 53.690 13.590 53.990 14.440 ;
        RECT 55.690 13.590 55.990 14.440 ;
        RECT 57.690 13.590 57.990 14.440 ;
        RECT 59.690 13.590 59.990 14.440 ;
        RECT 61.690 13.590 61.990 14.440 ;
        RECT 63.690 13.590 63.990 14.440 ;
        RECT 65.690 13.590 65.990 14.440 ;
        RECT 67.690 13.590 67.990 14.440 ;
        RECT 69.690 13.590 69.990 14.440 ;
        RECT 71.690 13.590 71.990 14.440 ;
        RECT 73.690 13.590 73.990 14.440 ;
        RECT 87.125 13.590 87.425 14.440 ;
        RECT 89.125 13.590 89.425 14.440 ;
        RECT 91.125 13.590 91.425 14.440 ;
        RECT 93.125 13.590 93.425 14.440 ;
        RECT 95.125 13.590 95.425 14.440 ;
        RECT 97.125 13.590 97.425 14.440 ;
        RECT 99.125 13.590 99.425 14.440 ;
        RECT 101.125 13.590 101.425 14.440 ;
        RECT 103.125 13.590 103.425 14.440 ;
        RECT 105.125 13.590 105.425 14.440 ;
        RECT 107.125 13.590 107.425 14.440 ;
        RECT 109.125 13.590 109.425 14.440 ;
        RECT 111.125 13.590 111.425 14.440 ;
        RECT 113.125 13.590 113.425 14.440 ;
        RECT 115.125 13.590 115.425 14.440 ;
        RECT 117.125 13.590 117.425 14.440 ;
        RECT 119.125 13.590 119.425 14.440 ;
        RECT 121.125 13.590 121.425 14.440 ;
        RECT 123.125 13.590 123.425 14.440 ;
        RECT 125.125 13.590 125.425 14.440 ;
        RECT 127.125 13.590 127.425 14.440 ;
        RECT 129.125 13.590 129.425 14.440 ;
        RECT 131.125 13.590 131.425 14.440 ;
        RECT 133.125 13.590 133.425 14.440 ;
        RECT 135.125 13.590 135.425 14.440 ;
        RECT 137.125 13.590 137.425 14.440 ;
        RECT 139.125 13.590 139.425 14.440 ;
        RECT 141.125 13.590 141.425 14.440 ;
        RECT 143.125 13.590 143.425 14.440 ;
        RECT 145.125 13.590 145.425 14.440 ;
        RECT 147.125 13.590 147.425 14.440 ;
        RECT 149.125 13.590 149.425 14.440 ;
        RECT 151.125 13.590 151.425 14.440 ;
        RECT 153.125 13.590 153.425 14.440 ;
        RECT 7.340 12.590 8.340 13.590 ;
        RECT 9.340 12.590 10.340 13.590 ;
        RECT 11.340 12.590 12.340 13.590 ;
        RECT 13.340 12.590 14.340 13.590 ;
        RECT 15.340 12.590 16.340 13.590 ;
        RECT 17.340 12.590 18.340 13.590 ;
        RECT 19.340 12.590 20.340 13.590 ;
        RECT 21.340 12.590 22.340 13.590 ;
        RECT 23.340 12.590 24.340 13.590 ;
        RECT 25.340 12.590 26.340 13.590 ;
        RECT 27.340 12.590 28.340 13.590 ;
        RECT 29.340 12.590 30.340 13.590 ;
        RECT 31.340 12.590 32.340 13.590 ;
        RECT 33.340 12.590 34.340 13.590 ;
        RECT 35.340 12.590 36.340 13.590 ;
        RECT 37.340 12.590 38.340 13.590 ;
        RECT 39.340 12.590 40.340 13.590 ;
        RECT 41.340 12.590 42.340 13.590 ;
        RECT 43.340 12.590 44.340 13.590 ;
        RECT 45.340 12.590 46.340 13.590 ;
        RECT 47.340 12.590 48.340 13.590 ;
        RECT 49.340 12.590 50.340 13.590 ;
        RECT 51.340 12.590 52.340 13.590 ;
        RECT 53.340 12.590 54.340 13.590 ;
        RECT 55.340 12.590 56.340 13.590 ;
        RECT 57.340 12.590 58.340 13.590 ;
        RECT 59.340 12.590 60.340 13.590 ;
        RECT 61.340 12.590 62.340 13.590 ;
        RECT 63.340 12.590 64.340 13.590 ;
        RECT 65.340 12.590 66.340 13.590 ;
        RECT 67.340 12.590 68.340 13.590 ;
        RECT 69.340 12.590 70.340 13.590 ;
        RECT 71.340 12.590 72.340 13.590 ;
        RECT 73.340 12.590 74.340 13.590 ;
        RECT 86.775 12.590 87.775 13.590 ;
        RECT 88.775 12.590 89.775 13.590 ;
        RECT 90.775 12.590 91.775 13.590 ;
        RECT 92.775 12.590 93.775 13.590 ;
        RECT 94.775 12.590 95.775 13.590 ;
        RECT 96.775 12.590 97.775 13.590 ;
        RECT 98.775 12.590 99.775 13.590 ;
        RECT 100.775 12.590 101.775 13.590 ;
        RECT 102.775 12.590 103.775 13.590 ;
        RECT 104.775 12.590 105.775 13.590 ;
        RECT 106.775 12.590 107.775 13.590 ;
        RECT 108.775 12.590 109.775 13.590 ;
        RECT 110.775 12.590 111.775 13.590 ;
        RECT 112.775 12.590 113.775 13.590 ;
        RECT 114.775 12.590 115.775 13.590 ;
        RECT 116.775 12.590 117.775 13.590 ;
        RECT 118.775 12.590 119.775 13.590 ;
        RECT 120.775 12.590 121.775 13.590 ;
        RECT 122.775 12.590 123.775 13.590 ;
        RECT 124.775 12.590 125.775 13.590 ;
        RECT 126.775 12.590 127.775 13.590 ;
        RECT 128.775 12.590 129.775 13.590 ;
        RECT 130.775 12.590 131.775 13.590 ;
        RECT 132.775 12.590 133.775 13.590 ;
        RECT 134.775 12.590 135.775 13.590 ;
        RECT 136.775 12.590 137.775 13.590 ;
        RECT 138.775 12.590 139.775 13.590 ;
        RECT 140.775 12.590 141.775 13.590 ;
        RECT 142.775 12.590 143.775 13.590 ;
        RECT 144.775 12.590 145.775 13.590 ;
        RECT 146.775 12.590 147.775 13.590 ;
        RECT 148.775 12.590 149.775 13.590 ;
        RECT 150.775 12.590 151.775 13.590 ;
        RECT 152.775 12.590 153.775 13.590 ;
        RECT 7.690 11.740 7.990 12.590 ;
        RECT 9.690 11.740 9.990 12.590 ;
        RECT 11.690 11.740 11.990 12.590 ;
        RECT 13.690 11.740 13.990 12.590 ;
        RECT 15.690 11.740 15.990 12.590 ;
        RECT 17.690 11.740 17.990 12.590 ;
        RECT 19.690 11.740 19.990 12.590 ;
        RECT 21.690 11.740 21.990 12.590 ;
        RECT 23.690 11.740 23.990 12.590 ;
        RECT 25.690 11.740 25.990 12.590 ;
        RECT 27.690 11.740 27.990 12.590 ;
        RECT 29.690 11.740 29.990 12.590 ;
        RECT 31.690 11.740 31.990 12.590 ;
        RECT 33.690 11.740 33.990 12.590 ;
        RECT 35.690 11.740 35.990 12.590 ;
        RECT 37.690 11.740 37.990 12.590 ;
        RECT 39.690 11.740 39.990 12.590 ;
        RECT 41.690 11.740 41.990 12.590 ;
        RECT 43.690 11.740 43.990 12.590 ;
        RECT 45.690 11.740 45.990 12.590 ;
        RECT 47.690 11.740 47.990 12.590 ;
        RECT 49.690 11.740 49.990 12.590 ;
        RECT 51.690 11.740 51.990 12.590 ;
        RECT 53.690 11.740 53.990 12.590 ;
        RECT 55.690 11.740 55.990 12.590 ;
        RECT 57.690 11.740 57.990 12.590 ;
        RECT 59.690 11.740 59.990 12.590 ;
        RECT 61.690 11.740 61.990 12.590 ;
        RECT 63.690 11.740 63.990 12.590 ;
        RECT 65.690 11.740 65.990 12.590 ;
        RECT 67.690 11.740 67.990 12.590 ;
        RECT 69.690 11.740 69.990 12.590 ;
        RECT 71.690 11.740 71.990 12.590 ;
        RECT 73.690 11.740 73.990 12.590 ;
        RECT 87.125 11.740 87.425 12.590 ;
        RECT 89.125 11.740 89.425 12.590 ;
        RECT 91.125 11.740 91.425 12.590 ;
        RECT 93.125 11.740 93.425 12.590 ;
        RECT 95.125 11.740 95.425 12.590 ;
        RECT 97.125 11.740 97.425 12.590 ;
        RECT 99.125 11.740 99.425 12.590 ;
        RECT 101.125 11.740 101.425 12.590 ;
        RECT 103.125 11.740 103.425 12.590 ;
        RECT 105.125 11.740 105.425 12.590 ;
        RECT 107.125 11.740 107.425 12.590 ;
        RECT 109.125 11.740 109.425 12.590 ;
        RECT 111.125 11.740 111.425 12.590 ;
        RECT 113.125 11.740 113.425 12.590 ;
        RECT 115.125 11.740 115.425 12.590 ;
        RECT 117.125 11.740 117.425 12.590 ;
        RECT 119.125 11.740 119.425 12.590 ;
        RECT 121.125 11.740 121.425 12.590 ;
        RECT 123.125 11.740 123.425 12.590 ;
        RECT 125.125 11.740 125.425 12.590 ;
        RECT 127.125 11.740 127.425 12.590 ;
        RECT 129.125 11.740 129.425 12.590 ;
        RECT 131.125 11.740 131.425 12.590 ;
        RECT 133.125 11.740 133.425 12.590 ;
        RECT 135.125 11.740 135.425 12.590 ;
        RECT 137.125 11.740 137.425 12.590 ;
        RECT 139.125 11.740 139.425 12.590 ;
        RECT 141.125 11.740 141.425 12.590 ;
        RECT 143.125 11.740 143.425 12.590 ;
        RECT 145.125 11.740 145.425 12.590 ;
        RECT 147.125 11.740 147.425 12.590 ;
        RECT 149.125 11.740 149.425 12.590 ;
        RECT 151.125 11.740 151.425 12.590 ;
        RECT 153.125 11.740 153.425 12.590 ;
        RECT 7.340 10.740 8.340 11.740 ;
        RECT 9.340 10.740 10.340 11.740 ;
        RECT 11.340 10.740 12.340 11.740 ;
        RECT 13.340 10.740 14.340 11.740 ;
        RECT 15.340 10.740 16.340 11.740 ;
        RECT 17.340 10.740 18.340 11.740 ;
        RECT 19.340 10.740 20.340 11.740 ;
        RECT 21.340 10.740 22.340 11.740 ;
        RECT 23.340 10.740 24.340 11.740 ;
        RECT 25.340 10.740 26.340 11.740 ;
        RECT 27.340 10.740 28.340 11.740 ;
        RECT 29.340 10.740 30.340 11.740 ;
        RECT 31.340 10.740 32.340 11.740 ;
        RECT 33.340 10.740 34.340 11.740 ;
        RECT 35.340 10.740 36.340 11.740 ;
        RECT 37.340 10.740 38.340 11.740 ;
        RECT 39.340 10.740 40.340 11.740 ;
        RECT 41.340 10.740 42.340 11.740 ;
        RECT 43.340 10.740 44.340 11.740 ;
        RECT 45.340 10.740 46.340 11.740 ;
        RECT 47.340 10.740 48.340 11.740 ;
        RECT 49.340 10.740 50.340 11.740 ;
        RECT 51.340 10.740 52.340 11.740 ;
        RECT 53.340 10.740 54.340 11.740 ;
        RECT 55.340 10.740 56.340 11.740 ;
        RECT 57.340 10.740 58.340 11.740 ;
        RECT 59.340 10.740 60.340 11.740 ;
        RECT 61.340 10.740 62.340 11.740 ;
        RECT 63.340 10.740 64.340 11.740 ;
        RECT 65.340 10.740 66.340 11.740 ;
        RECT 67.340 10.740 68.340 11.740 ;
        RECT 69.340 10.740 70.340 11.740 ;
        RECT 71.340 10.740 72.340 11.740 ;
        RECT 73.340 10.740 74.340 11.740 ;
        RECT 86.775 10.740 87.775 11.740 ;
        RECT 88.775 10.740 89.775 11.740 ;
        RECT 90.775 10.740 91.775 11.740 ;
        RECT 92.775 10.740 93.775 11.740 ;
        RECT 94.775 10.740 95.775 11.740 ;
        RECT 96.775 10.740 97.775 11.740 ;
        RECT 98.775 10.740 99.775 11.740 ;
        RECT 100.775 10.740 101.775 11.740 ;
        RECT 102.775 10.740 103.775 11.740 ;
        RECT 104.775 10.740 105.775 11.740 ;
        RECT 106.775 10.740 107.775 11.740 ;
        RECT 108.775 10.740 109.775 11.740 ;
        RECT 110.775 10.740 111.775 11.740 ;
        RECT 112.775 10.740 113.775 11.740 ;
        RECT 114.775 10.740 115.775 11.740 ;
        RECT 116.775 10.740 117.775 11.740 ;
        RECT 118.775 10.740 119.775 11.740 ;
        RECT 120.775 10.740 121.775 11.740 ;
        RECT 122.775 10.740 123.775 11.740 ;
        RECT 124.775 10.740 125.775 11.740 ;
        RECT 126.775 10.740 127.775 11.740 ;
        RECT 128.775 10.740 129.775 11.740 ;
        RECT 130.775 10.740 131.775 11.740 ;
        RECT 132.775 10.740 133.775 11.740 ;
        RECT 134.775 10.740 135.775 11.740 ;
        RECT 136.775 10.740 137.775 11.740 ;
        RECT 138.775 10.740 139.775 11.740 ;
        RECT 140.775 10.740 141.775 11.740 ;
        RECT 142.775 10.740 143.775 11.740 ;
        RECT 144.775 10.740 145.775 11.740 ;
        RECT 146.775 10.740 147.775 11.740 ;
        RECT 148.775 10.740 149.775 11.740 ;
        RECT 150.775 10.740 151.775 11.740 ;
        RECT 152.775 10.740 153.775 11.740 ;
        RECT 7.690 9.890 7.990 10.740 ;
        RECT 9.690 9.890 9.990 10.740 ;
        RECT 11.690 9.890 11.990 10.740 ;
        RECT 13.690 9.890 13.990 10.740 ;
        RECT 15.690 9.890 15.990 10.740 ;
        RECT 17.690 9.890 17.990 10.740 ;
        RECT 19.690 9.890 19.990 10.740 ;
        RECT 21.690 9.890 21.990 10.740 ;
        RECT 23.690 9.890 23.990 10.740 ;
        RECT 25.690 9.890 25.990 10.740 ;
        RECT 27.690 9.890 27.990 10.740 ;
        RECT 29.690 9.890 29.990 10.740 ;
        RECT 31.690 9.890 31.990 10.740 ;
        RECT 33.690 9.890 33.990 10.740 ;
        RECT 35.690 9.890 35.990 10.740 ;
        RECT 37.690 9.890 37.990 10.740 ;
        RECT 39.690 9.890 39.990 10.740 ;
        RECT 41.690 9.890 41.990 10.740 ;
        RECT 43.690 9.890 43.990 10.740 ;
        RECT 45.690 9.890 45.990 10.740 ;
        RECT 47.690 9.890 47.990 10.740 ;
        RECT 49.690 9.890 49.990 10.740 ;
        RECT 51.690 9.890 51.990 10.740 ;
        RECT 53.690 9.890 53.990 10.740 ;
        RECT 55.690 9.890 55.990 10.740 ;
        RECT 57.690 9.890 57.990 10.740 ;
        RECT 59.690 9.890 59.990 10.740 ;
        RECT 61.690 9.890 61.990 10.740 ;
        RECT 63.690 9.890 63.990 10.740 ;
        RECT 65.690 9.890 65.990 10.740 ;
        RECT 67.690 9.890 67.990 10.740 ;
        RECT 69.690 9.890 69.990 10.740 ;
        RECT 71.690 9.890 71.990 10.740 ;
        RECT 73.690 9.890 73.990 10.740 ;
        RECT 87.125 9.890 87.425 10.740 ;
        RECT 89.125 9.890 89.425 10.740 ;
        RECT 91.125 9.890 91.425 10.740 ;
        RECT 93.125 9.890 93.425 10.740 ;
        RECT 95.125 9.890 95.425 10.740 ;
        RECT 97.125 9.890 97.425 10.740 ;
        RECT 99.125 9.890 99.425 10.740 ;
        RECT 101.125 9.890 101.425 10.740 ;
        RECT 103.125 9.890 103.425 10.740 ;
        RECT 105.125 9.890 105.425 10.740 ;
        RECT 107.125 9.890 107.425 10.740 ;
        RECT 109.125 9.890 109.425 10.740 ;
        RECT 111.125 9.890 111.425 10.740 ;
        RECT 113.125 9.890 113.425 10.740 ;
        RECT 115.125 9.890 115.425 10.740 ;
        RECT 117.125 9.890 117.425 10.740 ;
        RECT 119.125 9.890 119.425 10.740 ;
        RECT 121.125 9.890 121.425 10.740 ;
        RECT 123.125 9.890 123.425 10.740 ;
        RECT 125.125 9.890 125.425 10.740 ;
        RECT 127.125 9.890 127.425 10.740 ;
        RECT 129.125 9.890 129.425 10.740 ;
        RECT 131.125 9.890 131.425 10.740 ;
        RECT 133.125 9.890 133.425 10.740 ;
        RECT 135.125 9.890 135.425 10.740 ;
        RECT 137.125 9.890 137.425 10.740 ;
        RECT 139.125 9.890 139.425 10.740 ;
        RECT 141.125 9.890 141.425 10.740 ;
        RECT 143.125 9.890 143.425 10.740 ;
        RECT 145.125 9.890 145.425 10.740 ;
        RECT 147.125 9.890 147.425 10.740 ;
        RECT 149.125 9.890 149.425 10.740 ;
        RECT 151.125 9.890 151.425 10.740 ;
        RECT 153.125 9.890 153.425 10.740 ;
        RECT 7.340 8.890 8.340 9.890 ;
        RECT 9.340 8.890 10.340 9.890 ;
        RECT 11.340 8.890 12.340 9.890 ;
        RECT 13.340 8.890 14.340 9.890 ;
        RECT 15.340 8.890 16.340 9.890 ;
        RECT 17.340 8.890 18.340 9.890 ;
        RECT 19.340 8.890 20.340 9.890 ;
        RECT 21.340 8.890 22.340 9.890 ;
        RECT 23.340 8.890 24.340 9.890 ;
        RECT 25.340 8.890 26.340 9.890 ;
        RECT 27.340 8.890 28.340 9.890 ;
        RECT 29.340 8.890 30.340 9.890 ;
        RECT 31.340 8.890 32.340 9.890 ;
        RECT 33.340 8.890 34.340 9.890 ;
        RECT 35.340 8.890 36.340 9.890 ;
        RECT 37.340 8.890 38.340 9.890 ;
        RECT 39.340 8.890 40.340 9.890 ;
        RECT 41.340 8.890 42.340 9.890 ;
        RECT 43.340 8.890 44.340 9.890 ;
        RECT 45.340 8.890 46.340 9.890 ;
        RECT 47.340 8.890 48.340 9.890 ;
        RECT 49.340 8.890 50.340 9.890 ;
        RECT 51.340 8.890 52.340 9.890 ;
        RECT 53.340 8.890 54.340 9.890 ;
        RECT 55.340 8.890 56.340 9.890 ;
        RECT 57.340 8.890 58.340 9.890 ;
        RECT 59.340 8.890 60.340 9.890 ;
        RECT 61.340 8.890 62.340 9.890 ;
        RECT 63.340 8.890 64.340 9.890 ;
        RECT 65.340 8.890 66.340 9.890 ;
        RECT 67.340 8.890 68.340 9.890 ;
        RECT 69.340 8.890 70.340 9.890 ;
        RECT 71.340 8.890 72.340 9.890 ;
        RECT 73.340 8.890 74.340 9.890 ;
        RECT 86.775 8.890 87.775 9.890 ;
        RECT 88.775 8.890 89.775 9.890 ;
        RECT 90.775 8.890 91.775 9.890 ;
        RECT 92.775 8.890 93.775 9.890 ;
        RECT 94.775 8.890 95.775 9.890 ;
        RECT 96.775 8.890 97.775 9.890 ;
        RECT 98.775 8.890 99.775 9.890 ;
        RECT 100.775 8.890 101.775 9.890 ;
        RECT 102.775 8.890 103.775 9.890 ;
        RECT 104.775 8.890 105.775 9.890 ;
        RECT 106.775 8.890 107.775 9.890 ;
        RECT 108.775 8.890 109.775 9.890 ;
        RECT 110.775 8.890 111.775 9.890 ;
        RECT 112.775 8.890 113.775 9.890 ;
        RECT 114.775 8.890 115.775 9.890 ;
        RECT 116.775 8.890 117.775 9.890 ;
        RECT 118.775 8.890 119.775 9.890 ;
        RECT 120.775 8.890 121.775 9.890 ;
        RECT 122.775 8.890 123.775 9.890 ;
        RECT 124.775 8.890 125.775 9.890 ;
        RECT 126.775 8.890 127.775 9.890 ;
        RECT 128.775 8.890 129.775 9.890 ;
        RECT 130.775 8.890 131.775 9.890 ;
        RECT 132.775 8.890 133.775 9.890 ;
        RECT 134.775 8.890 135.775 9.890 ;
        RECT 136.775 8.890 137.775 9.890 ;
        RECT 138.775 8.890 139.775 9.890 ;
        RECT 140.775 8.890 141.775 9.890 ;
        RECT 142.775 8.890 143.775 9.890 ;
        RECT 144.775 8.890 145.775 9.890 ;
        RECT 146.775 8.890 147.775 9.890 ;
        RECT 148.775 8.890 149.775 9.890 ;
        RECT 150.775 8.890 151.775 9.890 ;
        RECT 152.775 8.890 153.775 9.890 ;
        RECT 7.690 8.040 7.990 8.890 ;
        RECT 9.690 8.040 9.990 8.890 ;
        RECT 11.690 8.040 11.990 8.890 ;
        RECT 13.690 8.040 13.990 8.890 ;
        RECT 15.690 8.040 15.990 8.890 ;
        RECT 17.690 8.040 17.990 8.890 ;
        RECT 19.690 8.040 19.990 8.890 ;
        RECT 21.690 8.040 21.990 8.890 ;
        RECT 23.690 8.040 23.990 8.890 ;
        RECT 25.690 8.040 25.990 8.890 ;
        RECT 27.690 8.040 27.990 8.890 ;
        RECT 29.690 8.040 29.990 8.890 ;
        RECT 31.690 8.040 31.990 8.890 ;
        RECT 33.690 8.040 33.990 8.890 ;
        RECT 35.690 8.040 35.990 8.890 ;
        RECT 37.690 8.040 37.990 8.890 ;
        RECT 39.690 8.040 39.990 8.890 ;
        RECT 41.690 8.040 41.990 8.890 ;
        RECT 43.690 8.040 43.990 8.890 ;
        RECT 45.690 8.040 45.990 8.890 ;
        RECT 47.690 8.040 47.990 8.890 ;
        RECT 49.690 8.040 49.990 8.890 ;
        RECT 51.690 8.040 51.990 8.890 ;
        RECT 53.690 8.040 53.990 8.890 ;
        RECT 55.690 8.040 55.990 8.890 ;
        RECT 57.690 8.040 57.990 8.890 ;
        RECT 59.690 8.040 59.990 8.890 ;
        RECT 61.690 8.040 61.990 8.890 ;
        RECT 63.690 8.040 63.990 8.890 ;
        RECT 65.690 8.040 65.990 8.890 ;
        RECT 67.690 8.040 67.990 8.890 ;
        RECT 69.690 8.040 69.990 8.890 ;
        RECT 71.690 8.040 71.990 8.890 ;
        RECT 73.690 8.040 73.990 8.890 ;
        RECT 87.125 8.040 87.425 8.890 ;
        RECT 89.125 8.040 89.425 8.890 ;
        RECT 91.125 8.040 91.425 8.890 ;
        RECT 93.125 8.040 93.425 8.890 ;
        RECT 95.125 8.040 95.425 8.890 ;
        RECT 97.125 8.040 97.425 8.890 ;
        RECT 99.125 8.040 99.425 8.890 ;
        RECT 101.125 8.040 101.425 8.890 ;
        RECT 103.125 8.040 103.425 8.890 ;
        RECT 105.125 8.040 105.425 8.890 ;
        RECT 107.125 8.040 107.425 8.890 ;
        RECT 109.125 8.040 109.425 8.890 ;
        RECT 111.125 8.040 111.425 8.890 ;
        RECT 113.125 8.040 113.425 8.890 ;
        RECT 115.125 8.040 115.425 8.890 ;
        RECT 117.125 8.040 117.425 8.890 ;
        RECT 119.125 8.040 119.425 8.890 ;
        RECT 121.125 8.040 121.425 8.890 ;
        RECT 123.125 8.040 123.425 8.890 ;
        RECT 125.125 8.040 125.425 8.890 ;
        RECT 127.125 8.040 127.425 8.890 ;
        RECT 129.125 8.040 129.425 8.890 ;
        RECT 131.125 8.040 131.425 8.890 ;
        RECT 133.125 8.040 133.425 8.890 ;
        RECT 135.125 8.040 135.425 8.890 ;
        RECT 137.125 8.040 137.425 8.890 ;
        RECT 139.125 8.040 139.425 8.890 ;
        RECT 141.125 8.040 141.425 8.890 ;
        RECT 143.125 8.040 143.425 8.890 ;
        RECT 145.125 8.040 145.425 8.890 ;
        RECT 147.125 8.040 147.425 8.890 ;
        RECT 149.125 8.040 149.425 8.890 ;
        RECT 151.125 8.040 151.425 8.890 ;
        RECT 153.125 8.040 153.425 8.890 ;
        RECT 7.340 7.040 8.340 8.040 ;
        RECT 9.340 7.040 10.340 8.040 ;
        RECT 11.340 7.040 12.340 8.040 ;
        RECT 13.340 7.040 14.340 8.040 ;
        RECT 15.340 7.040 16.340 8.040 ;
        RECT 17.340 7.040 18.340 8.040 ;
        RECT 19.340 7.040 20.340 8.040 ;
        RECT 21.340 7.040 22.340 8.040 ;
        RECT 23.340 7.040 24.340 8.040 ;
        RECT 25.340 7.040 26.340 8.040 ;
        RECT 27.340 7.040 28.340 8.040 ;
        RECT 29.340 7.040 30.340 8.040 ;
        RECT 31.340 7.040 32.340 8.040 ;
        RECT 33.340 7.040 34.340 8.040 ;
        RECT 35.340 7.040 36.340 8.040 ;
        RECT 37.340 7.040 38.340 8.040 ;
        RECT 39.340 7.040 40.340 8.040 ;
        RECT 41.340 7.040 42.340 8.040 ;
        RECT 43.340 7.040 44.340 8.040 ;
        RECT 45.340 7.040 46.340 8.040 ;
        RECT 47.340 7.040 48.340 8.040 ;
        RECT 49.340 7.040 50.340 8.040 ;
        RECT 51.340 7.040 52.340 8.040 ;
        RECT 53.340 7.040 54.340 8.040 ;
        RECT 55.340 7.040 56.340 8.040 ;
        RECT 57.340 7.040 58.340 8.040 ;
        RECT 59.340 7.040 60.340 8.040 ;
        RECT 61.340 7.040 62.340 8.040 ;
        RECT 63.340 7.040 64.340 8.040 ;
        RECT 65.340 7.040 66.340 8.040 ;
        RECT 67.340 7.040 68.340 8.040 ;
        RECT 69.340 7.040 70.340 8.040 ;
        RECT 71.340 7.040 72.340 8.040 ;
        RECT 73.340 7.040 74.340 8.040 ;
        RECT 86.775 7.040 87.775 8.040 ;
        RECT 88.775 7.040 89.775 8.040 ;
        RECT 90.775 7.040 91.775 8.040 ;
        RECT 92.775 7.040 93.775 8.040 ;
        RECT 94.775 7.040 95.775 8.040 ;
        RECT 96.775 7.040 97.775 8.040 ;
        RECT 98.775 7.040 99.775 8.040 ;
        RECT 100.775 7.040 101.775 8.040 ;
        RECT 102.775 7.040 103.775 8.040 ;
        RECT 104.775 7.040 105.775 8.040 ;
        RECT 106.775 7.040 107.775 8.040 ;
        RECT 108.775 7.040 109.775 8.040 ;
        RECT 110.775 7.040 111.775 8.040 ;
        RECT 112.775 7.040 113.775 8.040 ;
        RECT 114.775 7.040 115.775 8.040 ;
        RECT 116.775 7.040 117.775 8.040 ;
        RECT 118.775 7.040 119.775 8.040 ;
        RECT 120.775 7.040 121.775 8.040 ;
        RECT 122.775 7.040 123.775 8.040 ;
        RECT 124.775 7.040 125.775 8.040 ;
        RECT 126.775 7.040 127.775 8.040 ;
        RECT 128.775 7.040 129.775 8.040 ;
        RECT 130.775 7.040 131.775 8.040 ;
        RECT 132.775 7.040 133.775 8.040 ;
        RECT 134.775 7.040 135.775 8.040 ;
        RECT 136.775 7.040 137.775 8.040 ;
        RECT 138.775 7.040 139.775 8.040 ;
        RECT 140.775 7.040 141.775 8.040 ;
        RECT 142.775 7.040 143.775 8.040 ;
        RECT 144.775 7.040 145.775 8.040 ;
        RECT 146.775 7.040 147.775 8.040 ;
        RECT 148.775 7.040 149.775 8.040 ;
        RECT 150.775 7.040 151.775 8.040 ;
        RECT 152.775 7.040 153.775 8.040 ;
        RECT 7.690 6.190 7.990 7.040 ;
        RECT 9.690 6.190 9.990 7.040 ;
        RECT 11.690 6.190 11.990 7.040 ;
        RECT 13.690 6.190 13.990 7.040 ;
        RECT 15.690 6.190 15.990 7.040 ;
        RECT 17.690 6.190 17.990 7.040 ;
        RECT 19.690 6.190 19.990 7.040 ;
        RECT 21.690 6.190 21.990 7.040 ;
        RECT 23.690 6.190 23.990 7.040 ;
        RECT 25.690 6.190 25.990 7.040 ;
        RECT 27.690 6.190 27.990 7.040 ;
        RECT 29.690 6.190 29.990 7.040 ;
        RECT 31.690 6.190 31.990 7.040 ;
        RECT 33.690 6.190 33.990 7.040 ;
        RECT 35.690 6.190 35.990 7.040 ;
        RECT 37.690 6.190 37.990 7.040 ;
        RECT 39.690 6.190 39.990 7.040 ;
        RECT 41.690 6.190 41.990 7.040 ;
        RECT 43.690 6.190 43.990 7.040 ;
        RECT 45.690 6.190 45.990 7.040 ;
        RECT 47.690 6.190 47.990 7.040 ;
        RECT 49.690 6.190 49.990 7.040 ;
        RECT 51.690 6.190 51.990 7.040 ;
        RECT 53.690 6.190 53.990 7.040 ;
        RECT 55.690 6.190 55.990 7.040 ;
        RECT 57.690 6.190 57.990 7.040 ;
        RECT 59.690 6.190 59.990 7.040 ;
        RECT 61.690 6.190 61.990 7.040 ;
        RECT 63.690 6.190 63.990 7.040 ;
        RECT 65.690 6.190 65.990 7.040 ;
        RECT 67.690 6.190 67.990 7.040 ;
        RECT 69.690 6.190 69.990 7.040 ;
        RECT 71.690 6.190 71.990 7.040 ;
        RECT 73.690 6.190 73.990 7.040 ;
        RECT 87.125 6.190 87.425 7.040 ;
        RECT 89.125 6.190 89.425 7.040 ;
        RECT 91.125 6.190 91.425 7.040 ;
        RECT 93.125 6.190 93.425 7.040 ;
        RECT 95.125 6.190 95.425 7.040 ;
        RECT 97.125 6.190 97.425 7.040 ;
        RECT 99.125 6.190 99.425 7.040 ;
        RECT 101.125 6.190 101.425 7.040 ;
        RECT 103.125 6.190 103.425 7.040 ;
        RECT 105.125 6.190 105.425 7.040 ;
        RECT 107.125 6.190 107.425 7.040 ;
        RECT 109.125 6.190 109.425 7.040 ;
        RECT 111.125 6.190 111.425 7.040 ;
        RECT 113.125 6.190 113.425 7.040 ;
        RECT 115.125 6.190 115.425 7.040 ;
        RECT 117.125 6.190 117.425 7.040 ;
        RECT 119.125 6.190 119.425 7.040 ;
        RECT 121.125 6.190 121.425 7.040 ;
        RECT 123.125 6.190 123.425 7.040 ;
        RECT 125.125 6.190 125.425 7.040 ;
        RECT 127.125 6.190 127.425 7.040 ;
        RECT 129.125 6.190 129.425 7.040 ;
        RECT 131.125 6.190 131.425 7.040 ;
        RECT 133.125 6.190 133.425 7.040 ;
        RECT 135.125 6.190 135.425 7.040 ;
        RECT 137.125 6.190 137.425 7.040 ;
        RECT 139.125 6.190 139.425 7.040 ;
        RECT 141.125 6.190 141.425 7.040 ;
        RECT 143.125 6.190 143.425 7.040 ;
        RECT 145.125 6.190 145.425 7.040 ;
        RECT 147.125 6.190 147.425 7.040 ;
        RECT 149.125 6.190 149.425 7.040 ;
        RECT 151.125 6.190 151.425 7.040 ;
        RECT 153.125 6.190 153.425 7.040 ;
        RECT 7.340 5.190 8.340 6.190 ;
        RECT 9.340 5.840 10.340 6.190 ;
        RECT 11.340 5.840 12.340 6.190 ;
        RECT 13.340 5.840 14.340 6.190 ;
        RECT 15.340 5.840 16.340 6.190 ;
        RECT 17.340 5.840 18.340 6.190 ;
        RECT 19.340 5.840 20.340 6.190 ;
        RECT 21.340 5.840 22.340 6.190 ;
        RECT 23.340 5.840 24.340 6.190 ;
        RECT 25.340 5.840 26.340 6.190 ;
        RECT 27.340 5.840 28.340 6.190 ;
        RECT 29.340 5.840 30.340 6.190 ;
        RECT 31.340 5.840 32.340 6.190 ;
        RECT 33.340 5.840 34.340 6.190 ;
        RECT 35.340 5.840 36.340 6.190 ;
        RECT 37.340 5.840 38.340 6.190 ;
        RECT 39.340 5.840 40.340 6.190 ;
        RECT 41.340 5.840 42.340 6.190 ;
        RECT 43.340 5.840 44.340 6.190 ;
        RECT 45.340 5.840 46.340 6.190 ;
        RECT 47.340 5.840 48.340 6.190 ;
        RECT 49.340 5.840 50.340 6.190 ;
        RECT 51.340 5.840 52.340 6.190 ;
        RECT 53.340 5.840 54.340 6.190 ;
        RECT 55.340 5.840 56.340 6.190 ;
        RECT 57.340 5.840 58.340 6.190 ;
        RECT 59.340 5.840 60.340 6.190 ;
        RECT 61.340 5.840 62.340 6.190 ;
        RECT 63.340 5.840 64.340 6.190 ;
        RECT 65.340 5.840 66.340 6.190 ;
        RECT 67.340 5.840 68.340 6.190 ;
        RECT 69.340 5.840 70.340 6.190 ;
        RECT 71.340 5.840 72.340 6.190 ;
        RECT 9.340 5.540 72.340 5.840 ;
        RECT 9.340 5.190 10.340 5.540 ;
        RECT 11.340 5.190 12.340 5.540 ;
        RECT 13.340 5.190 14.340 5.540 ;
        RECT 15.340 5.190 16.340 5.540 ;
        RECT 17.340 5.190 18.340 5.540 ;
        RECT 19.340 5.190 20.340 5.540 ;
        RECT 21.340 5.190 22.340 5.540 ;
        RECT 23.340 5.190 24.340 5.540 ;
        RECT 25.340 5.190 26.340 5.540 ;
        RECT 27.340 5.190 28.340 5.540 ;
        RECT 29.340 5.190 30.340 5.540 ;
        RECT 31.340 5.190 32.340 5.540 ;
        RECT 33.340 5.190 34.340 5.540 ;
        RECT 35.340 5.190 36.340 5.540 ;
        RECT 37.340 5.190 38.340 5.540 ;
        RECT 39.340 5.190 40.340 5.540 ;
        RECT 41.340 5.190 42.340 5.540 ;
        RECT 43.340 5.190 44.340 5.540 ;
        RECT 45.340 5.190 46.340 5.540 ;
        RECT 47.340 5.190 48.340 5.540 ;
        RECT 49.340 5.190 50.340 5.540 ;
        RECT 51.340 5.190 52.340 5.540 ;
        RECT 53.340 5.190 54.340 5.540 ;
        RECT 55.340 5.190 56.340 5.540 ;
        RECT 57.340 5.190 58.340 5.540 ;
        RECT 59.340 5.190 60.340 5.540 ;
        RECT 61.340 5.190 62.340 5.540 ;
        RECT 63.340 5.190 64.340 5.540 ;
        RECT 65.340 5.190 66.340 5.540 ;
        RECT 67.340 5.190 68.340 5.540 ;
        RECT 69.340 5.190 70.340 5.540 ;
        RECT 71.340 5.190 72.340 5.540 ;
        RECT 73.340 5.190 74.340 6.190 ;
        RECT 86.775 5.190 87.775 6.190 ;
        RECT 88.775 5.840 89.775 6.190 ;
        RECT 90.775 5.840 91.775 6.190 ;
        RECT 92.775 5.840 93.775 6.190 ;
        RECT 94.775 5.840 95.775 6.190 ;
        RECT 96.775 5.840 97.775 6.190 ;
        RECT 98.775 5.840 99.775 6.190 ;
        RECT 100.775 5.840 101.775 6.190 ;
        RECT 102.775 5.840 103.775 6.190 ;
        RECT 104.775 5.840 105.775 6.190 ;
        RECT 106.775 5.840 107.775 6.190 ;
        RECT 108.775 5.840 109.775 6.190 ;
        RECT 110.775 5.840 111.775 6.190 ;
        RECT 112.775 5.840 113.775 6.190 ;
        RECT 114.775 5.840 115.775 6.190 ;
        RECT 116.775 5.840 117.775 6.190 ;
        RECT 118.775 5.840 119.775 6.190 ;
        RECT 120.775 5.840 121.775 6.190 ;
        RECT 122.775 5.840 123.775 6.190 ;
        RECT 124.775 5.840 125.775 6.190 ;
        RECT 126.775 5.840 127.775 6.190 ;
        RECT 128.775 5.840 129.775 6.190 ;
        RECT 130.775 5.840 131.775 6.190 ;
        RECT 132.775 5.840 133.775 6.190 ;
        RECT 134.775 5.840 135.775 6.190 ;
        RECT 136.775 5.840 137.775 6.190 ;
        RECT 138.775 5.840 139.775 6.190 ;
        RECT 140.775 5.840 141.775 6.190 ;
        RECT 142.775 5.840 143.775 6.190 ;
        RECT 144.775 5.840 145.775 6.190 ;
        RECT 146.775 5.840 147.775 6.190 ;
        RECT 148.775 5.840 149.775 6.190 ;
        RECT 150.775 5.840 151.775 6.190 ;
        RECT 88.775 5.540 151.775 5.840 ;
        RECT 88.775 5.190 89.775 5.540 ;
        RECT 90.775 5.190 91.775 5.540 ;
        RECT 92.775 5.190 93.775 5.540 ;
        RECT 94.775 5.190 95.775 5.540 ;
        RECT 96.775 5.190 97.775 5.540 ;
        RECT 98.775 5.190 99.775 5.540 ;
        RECT 100.775 5.190 101.775 5.540 ;
        RECT 102.775 5.190 103.775 5.540 ;
        RECT 104.775 5.190 105.775 5.540 ;
        RECT 106.775 5.190 107.775 5.540 ;
        RECT 108.775 5.190 109.775 5.540 ;
        RECT 110.775 5.190 111.775 5.540 ;
        RECT 112.775 5.190 113.775 5.540 ;
        RECT 114.775 5.190 115.775 5.540 ;
        RECT 116.775 5.190 117.775 5.540 ;
        RECT 118.775 5.190 119.775 5.540 ;
        RECT 120.775 5.190 121.775 5.540 ;
        RECT 122.775 5.190 123.775 5.540 ;
        RECT 124.775 5.190 125.775 5.540 ;
        RECT 126.775 5.190 127.775 5.540 ;
        RECT 128.775 5.190 129.775 5.540 ;
        RECT 130.775 5.190 131.775 5.540 ;
        RECT 132.775 5.190 133.775 5.540 ;
        RECT 134.775 5.190 135.775 5.540 ;
        RECT 136.775 5.190 137.775 5.540 ;
        RECT 138.775 5.190 139.775 5.540 ;
        RECT 140.775 5.190 141.775 5.540 ;
        RECT 142.775 5.190 143.775 5.540 ;
        RECT 144.775 5.190 145.775 5.540 ;
        RECT 146.775 5.190 147.775 5.540 ;
        RECT 148.775 5.190 149.775 5.540 ;
        RECT 150.775 5.190 151.775 5.540 ;
        RECT 152.775 5.190 153.775 6.190 ;
        RECT 7.690 4.790 7.990 5.190 ;
        RECT 9.690 4.790 9.990 5.190 ;
        RECT 11.690 4.790 11.990 5.190 ;
        RECT 13.690 4.790 13.990 5.190 ;
        RECT 15.690 4.790 15.990 5.190 ;
        RECT 17.690 4.790 17.990 5.190 ;
        RECT 19.690 4.790 19.990 5.190 ;
        RECT 21.690 4.790 21.990 5.190 ;
        RECT 23.690 4.790 23.990 5.190 ;
        RECT 25.690 4.790 25.990 5.190 ;
        RECT 27.690 4.790 27.990 5.190 ;
        RECT 29.690 4.790 29.990 5.190 ;
        RECT 31.690 4.790 31.990 5.190 ;
        RECT 33.690 4.790 33.990 5.190 ;
        RECT 35.690 4.790 35.990 5.190 ;
        RECT 37.690 4.790 37.990 5.190 ;
        RECT 39.690 4.790 39.990 5.190 ;
        RECT 41.690 4.790 41.990 5.190 ;
        RECT 43.690 4.790 43.990 5.190 ;
        RECT 45.690 4.790 45.990 5.190 ;
        RECT 47.690 4.790 47.990 5.190 ;
        RECT 49.690 4.790 49.990 5.190 ;
        RECT 51.690 4.790 51.990 5.190 ;
        RECT 53.690 4.790 53.990 5.190 ;
        RECT 55.690 4.790 55.990 5.190 ;
        RECT 57.690 4.790 57.990 5.190 ;
        RECT 59.690 4.790 59.990 5.190 ;
        RECT 61.690 4.790 61.990 5.190 ;
        RECT 63.690 4.790 63.990 5.190 ;
        RECT 65.690 4.790 65.990 5.190 ;
        RECT 67.690 4.790 67.990 5.190 ;
        RECT 69.690 4.790 69.990 5.190 ;
        RECT 71.690 4.790 71.990 5.190 ;
        RECT 73.690 4.790 73.990 5.190 ;
        RECT 87.125 4.790 87.425 5.190 ;
        RECT 89.125 4.790 89.425 5.190 ;
        RECT 91.125 4.790 91.425 5.190 ;
        RECT 93.125 4.790 93.425 5.190 ;
        RECT 95.125 4.790 95.425 5.190 ;
        RECT 97.125 4.790 97.425 5.190 ;
        RECT 99.125 4.790 99.425 5.190 ;
        RECT 101.125 4.790 101.425 5.190 ;
        RECT 103.125 4.790 103.425 5.190 ;
        RECT 105.125 4.790 105.425 5.190 ;
        RECT 107.125 4.790 107.425 5.190 ;
        RECT 109.125 4.790 109.425 5.190 ;
        RECT 111.125 4.790 111.425 5.190 ;
        RECT 113.125 4.790 113.425 5.190 ;
        RECT 115.125 4.790 115.425 5.190 ;
        RECT 117.125 4.790 117.425 5.190 ;
        RECT 119.125 4.790 119.425 5.190 ;
        RECT 121.125 4.790 121.425 5.190 ;
        RECT 123.125 4.790 123.425 5.190 ;
        RECT 125.125 4.790 125.425 5.190 ;
        RECT 127.125 4.790 127.425 5.190 ;
        RECT 129.125 4.790 129.425 5.190 ;
        RECT 131.125 4.790 131.425 5.190 ;
        RECT 133.125 4.790 133.425 5.190 ;
        RECT 135.125 4.790 135.425 5.190 ;
        RECT 137.125 4.790 137.425 5.190 ;
        RECT 139.125 4.790 139.425 5.190 ;
        RECT 141.125 4.790 141.425 5.190 ;
        RECT 143.125 4.790 143.425 5.190 ;
        RECT 145.125 4.790 145.425 5.190 ;
        RECT 147.125 4.790 147.425 5.190 ;
        RECT 149.125 4.790 149.425 5.190 ;
        RECT 151.125 4.790 151.425 5.190 ;
        RECT 153.125 4.790 153.425 5.190 ;
        RECT 68.090 1.000 68.990 2.500 ;
        RECT 90.170 1.000 91.070 1.600 ;
        RECT 112.250 1.000 113.150 3.450 ;
        RECT 134.330 1.000 135.230 4.100 ;
        RECT 154.265 1.000 155.165 4.750 ;
        RECT 154.265 0.100 156.410 1.000 ;
  END
END tt_um_rnunes2311_12bit_sar_adc
END LIBRARY

