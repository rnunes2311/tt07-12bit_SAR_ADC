magic
tech sky130A
magscale 1 2
timestamp 1715420247
<< metal2 >>
rect 2970 44685 3030 44695
rect 2970 44615 3030 44625
rect 2974 43952 3030 44615
rect 26890 44680 26950 44690
rect 26890 44610 26950 44620
rect 5362 44555 5422 44565
rect 5362 44485 5422 44495
rect 5366 43892 5422 44485
rect 24500 44450 24560 44460
rect 7754 44435 7814 44445
rect 24500 44380 24560 44390
rect 7754 44365 7814 44375
rect 7758 43892 7814 44365
rect 10146 44315 10208 44325
rect 19720 44320 19780 44330
rect 10206 44255 10208 44315
rect 10146 44245 10208 44255
rect 10150 43951 10208 44245
rect 19718 44260 19720 44318
rect 19718 44250 19780 44260
rect 12538 44195 12598 44205
rect 12538 44125 12598 44135
rect 12542 43972 12598 44125
rect 14930 44075 14990 44085
rect 14930 44005 14990 44015
rect 14934 43932 14990 44005
rect 17322 43960 17382 43970
rect 19718 43902 19774 44250
rect 22110 44190 22170 44200
rect 22108 44130 22110 44189
rect 22108 44120 22170 44130
rect 22108 43941 22166 44120
rect 17322 43890 17382 43900
rect 17326 43885 17382 43890
rect 24502 43702 24558 44380
rect 26894 43772 26950 44610
rect 29280 44570 29340 44580
rect 29340 44510 29342 44550
rect 29280 44500 29342 44510
rect 29286 43782 29342 44500
<< via2 >>
rect 2970 44625 3030 44685
rect 26890 44620 26950 44680
rect 5362 44495 5422 44555
rect 7754 44375 7814 44435
rect 24500 44390 24560 44450
rect 10146 44255 10206 44315
rect 19720 44260 19780 44320
rect 12538 44135 12598 44195
rect 14930 44015 14990 44075
rect 17322 43900 17382 43960
rect 22110 44130 22170 44190
rect 29280 44510 29340 44570
<< metal3 >>
rect 780 44750 790 44830
rect 870 44820 880 44830
rect 1510 44820 1520 44830
rect 870 44760 1520 44820
rect 870 44750 880 44760
rect 1510 44750 1520 44760
rect 1600 44820 1610 44830
rect 2250 44820 2260 44830
rect 1600 44760 2260 44820
rect 1600 44750 1610 44760
rect 2250 44750 2260 44760
rect 2340 44820 2350 44830
rect 2980 44820 2990 44830
rect 2340 44760 2990 44820
rect 2340 44750 2350 44760
rect 2980 44750 2990 44760
rect 3070 44820 3080 44830
rect 3720 44820 3730 44830
rect 3070 44760 3730 44820
rect 3070 44750 3080 44760
rect 3720 44750 3730 44760
rect 3810 44820 3820 44830
rect 4460 44820 4470 44830
rect 3810 44760 4470 44820
rect 3810 44750 3820 44760
rect 4460 44750 4470 44760
rect 4550 44820 4560 44830
rect 5190 44820 5200 44830
rect 4550 44760 5200 44820
rect 4550 44750 4560 44760
rect 5190 44750 5200 44760
rect 5280 44820 5290 44830
rect 5930 44820 5940 44830
rect 5280 44760 5940 44820
rect 5280 44750 5290 44760
rect 5930 44750 5940 44760
rect 6020 44820 6030 44830
rect 6670 44820 6680 44830
rect 6020 44760 6680 44820
rect 6020 44750 6030 44760
rect 6670 44750 6680 44760
rect 6760 44820 6770 44830
rect 7400 44820 7410 44830
rect 6760 44760 7410 44820
rect 6760 44750 6770 44760
rect 7400 44750 7410 44760
rect 7490 44820 7500 44830
rect 8140 44820 8150 44830
rect 7490 44760 8150 44820
rect 7490 44750 7500 44760
rect 8140 44750 8150 44760
rect 8230 44820 8240 44830
rect 8880 44820 8890 44830
rect 8230 44760 8890 44820
rect 8230 44750 8240 44760
rect 8880 44750 8890 44760
rect 8970 44820 8980 44830
rect 9610 44820 9620 44830
rect 8970 44760 9620 44820
rect 8970 44750 8980 44760
rect 9610 44750 9620 44760
rect 9700 44820 9710 44830
rect 10340 44820 10350 44830
rect 9700 44760 10350 44820
rect 9700 44750 9710 44760
rect 10340 44750 10350 44760
rect 10430 44820 10440 44830
rect 11080 44820 11090 44830
rect 10430 44760 11090 44820
rect 10430 44750 10440 44760
rect 11080 44750 11090 44760
rect 11170 44820 11180 44830
rect 11820 44820 11830 44830
rect 11170 44760 11830 44820
rect 11170 44750 11180 44760
rect 11820 44750 11830 44760
rect 11910 44820 11920 44830
rect 11910 44760 31840 44820
rect 11910 44750 11920 44760
rect 31830 44740 31840 44760
rect 31920 44740 31930 44820
rect 2960 44685 3040 44690
rect 2960 44625 2970 44685
rect 3030 44680 3040 44685
rect 13280 44680 13290 44700
rect 3030 44625 13290 44680
rect 2960 44620 13290 44625
rect 13370 44620 13380 44700
rect 26880 44680 26960 44685
rect 28004 44680 28014 44700
rect 26880 44620 26890 44680
rect 26950 44620 28014 44680
rect 28094 44620 28104 44700
rect 26880 44615 26960 44620
rect 14020 44560 14030 44580
rect 5352 44555 14030 44560
rect 5352 44495 5362 44555
rect 5422 44500 14030 44555
rect 14110 44500 14120 44580
rect 28740 44500 28750 44580
rect 28830 44560 28840 44580
rect 29270 44570 29350 44575
rect 29270 44560 29280 44570
rect 28830 44510 29280 44560
rect 29340 44510 29350 44570
rect 28830 44500 29350 44510
rect 5422 44495 5432 44500
rect 5352 44490 5432 44495
rect 14750 44440 14760 44460
rect 7744 44435 14760 44440
rect 7744 44375 7754 44435
rect 7814 44380 14760 44435
rect 14840 44380 14850 44460
rect 24490 44450 24570 44460
rect 24490 44390 24500 44450
rect 24560 44440 24570 44450
rect 29476 44440 29486 44460
rect 24560 44390 29486 44440
rect 24490 44380 29486 44390
rect 29566 44380 29576 44460
rect 7814 44375 7824 44380
rect 7744 44370 7824 44375
rect 15500 44320 15510 44340
rect 10136 44315 15510 44320
rect 10136 44255 10146 44315
rect 10206 44260 15510 44315
rect 15590 44260 15600 44340
rect 19710 44320 19790 44325
rect 30212 44320 30222 44340
rect 19710 44260 19720 44320
rect 19780 44260 30222 44320
rect 30302 44260 30312 44340
rect 10206 44255 10216 44260
rect 19710 44255 19790 44260
rect 10136 44250 10216 44255
rect 16230 44200 16240 44220
rect 12528 44195 16240 44200
rect 12528 44135 12538 44195
rect 12598 44140 16240 44195
rect 16320 44140 16330 44220
rect 30948 44200 30958 44220
rect 22100 44190 30958 44200
rect 12598 44135 12608 44140
rect 12528 44130 12608 44135
rect 22100 44130 22110 44190
rect 22170 44140 30958 44190
rect 31038 44140 31048 44220
rect 22170 44130 22180 44140
rect 22100 44125 22180 44130
rect 16960 44080 16970 44100
rect 14920 44075 16970 44080
rect 14920 44015 14930 44075
rect 14990 44020 16970 44075
rect 17050 44020 17060 44100
rect 14990 44015 15000 44020
rect 14920 44010 15000 44015
rect 17312 43960 17392 43965
rect 17700 43960 17710 43980
rect 17312 43900 17322 43960
rect 17382 43900 17710 43960
rect 17790 43900 17800 43980
rect 17312 43895 17392 43900
rect 658 440 718 860
rect 30833 830 30855 890
rect 30845 820 30855 830
rect 30925 820 30955 890
rect 31025 830 31055 890
rect 31025 820 31035 830
rect 26846 700 26868 760
rect 26858 690 26868 700
rect 26938 690 26968 760
rect 27038 700 27068 760
rect 27038 690 27048 700
rect 22430 570 22452 630
rect 22442 560 22452 570
rect 22522 560 22552 630
rect 22622 570 22652 630
rect 22622 560 22632 570
rect 658 380 13620 440
rect 13610 370 13620 380
rect 13690 370 13720 440
rect 13790 380 31370 440
rect 13790 370 13800 380
rect 31505 310 31565 790
rect 800 250 18036 310
rect 18026 240 18036 250
rect 18106 240 18136 310
rect 18206 250 31565 310
rect 18206 240 18216 250
<< via3 >>
rect 790 44750 870 44830
rect 1520 44750 1600 44830
rect 2260 44750 2340 44830
rect 2990 44750 3070 44830
rect 3730 44750 3810 44830
rect 4470 44750 4550 44830
rect 5200 44750 5280 44830
rect 5940 44750 6020 44830
rect 6680 44750 6760 44830
rect 7410 44750 7490 44830
rect 8150 44750 8230 44830
rect 8890 44750 8970 44830
rect 9620 44750 9700 44830
rect 10350 44750 10430 44830
rect 11090 44750 11170 44830
rect 11830 44750 11910 44830
rect 31840 44740 31920 44820
rect 13290 44620 13370 44700
rect 28014 44620 28094 44700
rect 14030 44500 14110 44580
rect 28750 44500 28830 44580
rect 14760 44380 14840 44460
rect 29486 44380 29566 44460
rect 15510 44260 15590 44340
rect 30222 44260 30302 44340
rect 16240 44140 16320 44220
rect 30958 44140 31038 44220
rect 16970 44020 17050 44100
rect 17710 43900 17790 43980
rect 30855 820 30925 890
rect 30955 820 31025 890
rect 26868 690 26938 760
rect 26968 690 27038 760
rect 22452 560 22522 630
rect 22552 560 22622 630
rect 13620 370 13690 440
rect 13720 370 13790 440
rect 18036 240 18106 310
rect 18136 240 18206 310
<< metal4 >>
rect 798 44831 858 45152
rect 1534 44831 1594 45152
rect 2270 44831 2330 45152
rect 3006 44831 3066 45152
rect 3742 44831 3802 45152
rect 4478 44831 4538 45152
rect 5214 44831 5274 45152
rect 5950 44831 6010 45152
rect 6686 44831 6746 45152
rect 7422 44831 7482 45152
rect 8158 44831 8218 45152
rect 8894 44831 8954 45152
rect 9630 44831 9690 45152
rect 10366 44831 10426 45152
rect 11102 44831 11162 45152
rect 11838 44831 11898 45152
rect 12574 44952 12634 45152
rect 789 44830 871 44831
rect 789 44750 790 44830
rect 870 44750 871 44830
rect 789 44749 871 44750
rect 1519 44830 1601 44831
rect 1519 44750 1520 44830
rect 1600 44750 1601 44830
rect 1519 44749 1601 44750
rect 2259 44830 2341 44831
rect 2259 44750 2260 44830
rect 2340 44750 2341 44830
rect 2259 44749 2341 44750
rect 2989 44830 3071 44831
rect 2989 44750 2990 44830
rect 3070 44750 3071 44830
rect 2989 44749 3071 44750
rect 3729 44830 3811 44831
rect 3729 44750 3730 44830
rect 3810 44750 3811 44830
rect 3729 44749 3811 44750
rect 4469 44830 4551 44831
rect 4469 44750 4470 44830
rect 4550 44750 4551 44830
rect 4469 44749 4551 44750
rect 5199 44830 5281 44831
rect 5199 44750 5200 44830
rect 5280 44750 5281 44830
rect 5199 44749 5281 44750
rect 5939 44830 6021 44831
rect 5939 44750 5940 44830
rect 6020 44750 6021 44830
rect 5939 44749 6021 44750
rect 6679 44830 6761 44831
rect 6679 44750 6680 44830
rect 6760 44750 6761 44830
rect 6679 44749 6761 44750
rect 7409 44830 7491 44831
rect 7409 44750 7410 44830
rect 7490 44750 7491 44830
rect 7409 44749 7491 44750
rect 8149 44830 8231 44831
rect 8149 44750 8150 44830
rect 8230 44750 8231 44830
rect 8149 44749 8231 44750
rect 8889 44830 8971 44831
rect 8889 44750 8890 44830
rect 8970 44750 8971 44830
rect 8889 44749 8971 44750
rect 9619 44830 9701 44831
rect 9619 44750 9620 44830
rect 9700 44750 9701 44830
rect 9619 44749 9701 44750
rect 10349 44830 10431 44831
rect 10349 44750 10350 44830
rect 10430 44750 10431 44830
rect 10349 44749 10431 44750
rect 11089 44830 11171 44831
rect 11089 44750 11090 44830
rect 11170 44750 11171 44830
rect 11089 44749 11171 44750
rect 11829 44830 11911 44831
rect 11829 44750 11830 44830
rect 11910 44750 11911 44830
rect 11829 44749 11911 44750
rect 13310 44701 13370 45152
rect 13289 44700 13371 44701
rect 13289 44620 13290 44700
rect 13370 44620 13371 44700
rect 13289 44619 13371 44620
rect 14046 44581 14106 45152
rect 14029 44580 14111 44581
rect 14029 44500 14030 44580
rect 14110 44500 14111 44580
rect 14029 44499 14111 44500
rect 14782 44461 14842 45152
rect 14759 44460 14842 44461
rect 14759 44380 14760 44460
rect 14840 44430 14842 44460
rect 14840 44380 14841 44430
rect 14759 44379 14841 44380
rect 15518 44341 15578 45152
rect 15509 44340 15591 44341
rect 15509 44260 15510 44340
rect 15590 44260 15591 44340
rect 15509 44259 15591 44260
rect 16254 44221 16314 45152
rect 16239 44220 16321 44221
rect 200 43030 500 44152
rect 16239 44140 16240 44220
rect 16320 44140 16321 44220
rect 16239 44139 16321 44140
rect 16990 44101 17050 45152
rect 16969 44100 17051 44101
rect 16969 44020 16970 44100
rect 17050 44020 17051 44100
rect 16969 44019 17051 44020
rect 17726 43981 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44701 28090 45152
rect 28013 44700 28095 44701
rect 28013 44620 28014 44700
rect 28094 44620 28095 44700
rect 28013 44619 28095 44620
rect 28766 44581 28826 45152
rect 28749 44580 28831 44581
rect 28749 44500 28750 44580
rect 28830 44500 28831 44580
rect 28749 44499 28831 44500
rect 29502 44461 29562 45152
rect 29485 44460 29567 44461
rect 29485 44380 29486 44460
rect 29566 44380 29567 44460
rect 29485 44379 29567 44380
rect 30238 44341 30298 45152
rect 30221 44340 30303 44341
rect 30221 44260 30222 44340
rect 30302 44260 30303 44340
rect 30221 44259 30303 44260
rect 30974 44221 31034 45152
rect 31710 44952 31770 45152
rect 31700 44820 32000 44830
rect 31700 44740 31840 44820
rect 31920 44740 32000 44820
rect 30957 44220 31039 44221
rect 30957 44140 30958 44220
rect 31038 44140 31039 44220
rect 30957 44139 31039 44140
rect 17709 43980 17791 43981
rect 17709 43900 17710 43980
rect 17790 43900 17791 43980
rect 17709 43899 17791 43900
rect 31700 43046 32000 44740
rect 200 42730 6090 43030
rect 6615 42746 32000 43046
rect 200 41080 500 42730
rect 200 40780 6120 41080
rect 200 39090 500 40780
rect 200 38790 6040 39090
rect 200 36910 500 38790
rect 31700 38296 32000 42746
rect 6625 37996 32000 38296
rect 5867 36910 5891 36954
rect 200 36610 6070 36910
rect 31700 36806 32000 37996
rect 200 34450 500 36610
rect 28699 36506 32000 36806
rect 200 34150 6110 34450
rect 200 31890 500 34150
rect 31700 33533 32000 36506
rect 28663 33233 32000 33533
rect 29008 33188 29009 33233
rect 200 31590 6100 31890
rect 200 1000 500 31590
rect 31700 1000 32000 33233
rect 30853 890 31033 902
rect 30853 820 30855 890
rect 30925 820 30955 890
rect 31025 820 31033 890
rect 26866 760 27046 772
rect 26866 690 26868 760
rect 26938 690 26968 760
rect 27038 690 27046 760
rect 22450 630 22630 642
rect 22450 560 22452 630
rect 22522 560 22552 630
rect 22622 560 22630 630
rect 13618 440 13798 450
rect 13618 370 13620 440
rect 13690 370 13720 440
rect 13790 370 13798 440
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 370
rect 18034 310 18214 320
rect 18034 240 18036 310
rect 18106 240 18136 310
rect 18206 240 18214 310
rect 18034 0 18214 240
rect 22450 0 22630 560
rect 26866 0 27046 690
rect 30853 200 31033 820
rect 30853 20 31462 200
rect 31282 0 31462 20
use SAR_ADC_12bit/layout/SAR_ADC_12bit  SAR_ADC_12bit_0 SAR_ADC_12bit/layout
timestamp 1715420247
transform 1 0 5968 0 1 -4142
box -5320 4712 25607 48195
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 31700 1000 32000 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
